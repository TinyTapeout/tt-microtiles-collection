/* Automatically generated from https://wokwi.com/projects/395357890431011841 */

`default_nettype none

module tt_um_wokwi_395357890431011841(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = ui_in[1];
  wire net3 = ui_in[2];
  wire net4;
  wire net5;
  wire net6;
  wire net7;
  wire net8;
  wire net9;
  wire net10;
  wire net11;
  wire net12 = 1'b0;
  wire net13 = 1'b1;
  wire net14 = 1'b1;
  wire net15 = 1'b0;
  wire net16 = 1'b1;
  wire net17;
  wire net18;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291;
  wire net292;
  wire net293;
  wire net294;
  wire net295;
  wire net296;
  wire net297;
  wire net298;
  wire net299;
  wire net300;
  wire net301;
  wire net302;
  wire net303;
  wire net304;
  wire net305;
  wire net306;
  wire net307;
  wire net308;
  wire net309;
  wire net310;
  wire net311;
  wire net312;
  wire net313;
  wire net314;
  wire net315;
  wire net316;
  wire net317;
  wire net318;
  wire net319;
  wire net320;
  wire net321;
  wire net322;
  wire net323;
  wire net324;
  wire net325;
  wire net326;
  wire net327;
  wire net328;
  wire net329;
  wire net330;
  wire net331;
  wire net332;
  wire net333;
  wire net334;
  wire net335;
  wire net336;
  wire net337;
  wire net338;
  wire net339;
  wire net340;
  wire net341;
  wire net342;
  wire net343;
  wire net344;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349;
  wire net350;
  wire net351;
  wire net352;
  wire net353;
  wire net354;
  wire net355;
  wire net356;
  wire net357;
  wire net358;
  wire net359;
  wire net360;
  wire net361;
  wire net362;
  wire net363;
  wire net364;
  wire net365;
  wire net366;
  wire net367;
  wire net368;
  wire net369;
  wire net370;
  wire net371;
  wire net372;
  wire net373;
  wire net374;
  wire net375;
  wire net376;
  wire net377;
  wire net378;
  wire net379;
  wire net380;
  wire net381;
  wire net382;
  wire net383;
  wire net384;
  wire net385;
  wire net386;
  wire net387;
  wire net388;
  wire net389;
  wire net390;
  wire net391;
  wire net392;
  wire net393;
  wire net394;
  wire net395;
  wire net396;
  wire net397;
  wire net398;
  wire net399;
  wire net400;
  wire net401;
  wire net402;
  wire net403;
  wire net404;
  wire net405;
  wire net406;
  wire net407;
  wire net408;
  wire net409;
  wire net410;
  wire net411;
  wire net412;
  wire net413;
  wire net414;
  wire net415;
  wire net416;
  wire net417;
  wire net418;
  wire net419;
  wire net420;
  wire net421;
  wire net422;
  wire net423;
  wire net424;
  wire net425;
  wire net426;
  wire net427;
  wire net428;
  wire net429;
  wire net430;
  wire net431;
  wire net432;
  wire net433;
  wire net434;
  wire net435;
  wire net436;
  wire net437;
  wire net438;
  wire net439;
  wire net440;
  wire net441;
  wire net442;
  wire net443;
  wire net444;
  wire net445;
  wire net446;
  wire net447;
  wire net448;
  wire net449;
  wire net450;
  wire net451;
  wire net452;
  wire net453;
  wire net454;
  wire net455;
  wire net456;
  wire net457;
  wire net458;
  wire net459;
  wire net460;
  wire net461;
  wire net462;
  wire net463;
  wire net464;
  wire net465;
  wire net466;
  wire net467;
  wire net468;
  wire net469;
  wire net470;
  wire net471;
  wire net472;
  wire net473;
  wire net474;
  wire net475;
  wire net476;
  wire net477;
  wire net478;
  wire net479;
  wire net480;
  wire net481;
  wire net482;
  wire net483;
  wire net484;
  wire net485;
  wire net486;
  wire net487;
  wire net488;
  wire net489;
  wire net490;
  wire net491;
  wire net492;
  wire net493;
  wire net494;
  wire net495;
  wire net496;
  wire net497;
  wire net498;
  wire net499;
  wire net500;
  wire net501;
  wire net502;
  wire net503;
  wire net504;
  wire net505;
  wire net506;
  wire net507;
  wire net508;
  wire net509;
  wire net510;
  wire net511;
  wire net512;
  wire net513;
  wire net514;
  wire net515;
  wire net516;
  wire net517;
  wire net518;
  wire net519;
  wire net520;
  wire net521;
  wire net522;
  wire net523;
  wire net524;
  wire net525;
  wire net526;
  wire net527;
  wire net528;
  wire net529;
  wire net530;
  wire net531;
  wire net532;
  wire net533;
  wire net534;
  wire net535;
  wire net536;
  wire net537;
  wire net538;
  wire net539;
  wire net540;
  wire net541;
  wire net542;
  wire net543;
  wire net544;
  wire net545;
  wire net546;
  wire net547;
  wire net548;
  wire net549;
  wire net550;
  wire net551;
  wire net552;
  wire net553;
  wire net554;
  wire net555;
  wire net556;
  wire net557;
  wire net558;
  wire net559;
  wire net560;
  wire net561;
  wire net562;
  wire net563;
  wire net564;
  wire net565;
  wire net566;
  wire net567;
  wire net568;
  wire net569;
  wire net570;
  wire net571;
  wire net572;
  wire net573;
  wire net574;
  wire net575;
  wire net576;
  wire net577;
  wire net578;
  wire net579;
  wire net580;
  wire net581;
  wire net582;
  wire net583;
  wire net584;
  wire net585;
  wire net586;
  wire net587;
  wire net588;
  wire net589;
  wire net590;
  wire net591;
  wire net592;
  wire net593;
  wire net594;
  wire net595;
  wire net596;
  wire net597;
  wire net598;
  wire net599;
  wire net600;
  wire net601;
  wire net602;
  wire net603;
  wire net604;
  wire net605;
  wire net606;
  wire net607;
  wire net608;
  wire net609;
  wire net610;
  wire net611;
  wire net612;
  wire net613;
  wire net614;
  wire net615;
  wire net616;
  wire net617;
  wire net618;
  wire net619;
  wire net620;
  wire net621;
  wire net622;
  wire net623;
  wire net624;
  wire net625;
  wire net626;
  wire net627;
  wire net628;
  wire net629;
  wire net630;
  wire net631;
  wire net632;
  wire net633;
  wire net634;
  wire net635;
  wire net636;
  wire net637;
  wire net638;
  wire net639;
  wire net640;
  wire net641;
  wire net642;
  wire net643;
  wire net644;
  wire net645;
  wire net646;
  wire net647;
  wire net648;
  wire net649;
  wire net650;
  wire net651;
  wire net652;
  wire net653;
  wire net654;
  wire net655;
  wire net656;
  wire net657;
  wire net658;
  wire net659;
  wire net660;
  wire net661;
  wire net662;
  wire net663;
  wire net664;
  wire net665;
  wire net666;
  wire net667;
  wire net668;
  wire net669;
  wire net670;
  wire net671;
  wire net672;
  wire net673;
  wire net674;
  wire net675;
  wire net676;
  wire net677;
  wire net678;
  wire net679;
  wire net680;
  wire net681;
  wire net682;
  wire net683;
  wire net684;
  wire net685;
  wire net686;
  wire net687;
  wire net688;
  wire net689;
  wire net690;
  wire net691;
  wire net692;
  wire net693;
  wire net694;
  wire net695;
  wire net696;
  wire net697;
  wire net698;
  wire net699;
  wire net700;
  wire net701;
  wire net702;
  wire net703;
  wire net704;
  wire net705;
  wire net706;
  wire net707;
  wire net708;
  wire net709;
  wire net710;
  wire net711;
  wire net712;
  wire net713;
  wire net714;
  wire net715;
  wire net716;
  wire net717;
  wire net718;
  wire net719;
  wire net720;
  wire net721;
  wire net722;
  wire net723;
  wire net724;
  wire net725;
  wire net726;
  wire net727;
  wire net728;
  wire net729;
  wire net730;
  wire net731;
  wire net732;
  wire net733;
  wire net734;
  wire net735;
  wire net736;
  wire net737;
  wire net738;
  wire net739;
  wire net740;
  wire net741;
  wire net742;
  wire net743;
  wire net744;
  wire net745;
  wire net746;
  wire net747;
  wire net748;
  wire net749;
  wire net750;
  wire net751;
  wire net752;
  wire net753;
  wire net754;
  wire net755;
  wire net756;
  wire net757;
  wire net758;
  wire net759;
  wire net760;
  wire net761;
  wire net762;
  wire net763;
  wire net764;
  wire net765;
  wire net766;
  wire net767;
  wire net768;
  wire net769;
  wire net770;
  wire net771;
  wire net772;
  wire net773;
  wire net774;
  wire net775;
  wire net776;
  wire net777;
  wire net778;
  wire net779;
  wire net780;
  wire net781;
  wire net782;
  wire net783;
  wire net784;
  wire net785;
  wire net786;
  wire net787;
  wire net788;
  wire net789;
  wire net790;
  wire net791;
  wire net792;
  wire net793;
  wire net794;
  wire net795;
  wire net796;
  wire net797;
  wire net798;
  wire net799;
  wire net800;
  wire net801;
  wire net802;
  wire net803;
  wire net804;
  wire net805;
  wire net806;
  wire net807;
  wire net808;
  wire net809;
  wire net810;
  wire net811;
  wire net812;
  wire net813;
  wire net814;
  wire net815;
  wire net816;
  wire net817;
  wire net818;
  wire net819;
  wire net820;
  wire net821;
  wire net822;
  wire net823;
  wire net824;
  wire net825;
  wire net826;
  wire net827;
  wire net828;
  wire net829;
  wire net830;
  wire net831;
  wire net832;
  wire net833;
  wire net834;
  wire net835;
  wire net836;
  wire net837;
  wire net838;
  wire net839;
  wire net840;
  wire net841;
  wire net842;
  wire net843;
  wire net844;
  wire net845;
  wire net846;
  wire net847;
  wire net848;
  wire net849;
  wire net850;
  wire net851;
  wire net852;
  wire net853;
  wire net854;
  wire net855;
  wire net856;
  wire net857;
  wire net858;
  wire net859;
  wire net860;
  wire net861;
  wire net862;
  wire net863;
  wire net864;
  wire net865;
  wire net866;
  wire net867;
  wire net868;
  wire net869;
  wire net870;
  wire net871;
  wire net872;
  wire net873;
  wire net874;
  wire net875;
  wire net876;
  wire net877;
  wire net878;
  wire net879;
  wire net880;
  wire net881;
  wire net882;
  wire net883;
  wire net884;
  wire net885;
  wire net886;
  wire net887;
  wire net888;
  wire net889;

  assign uo_out[0] = net4;
  assign uo_out[1] = net5;
  assign uo_out[2] = net6;
  assign uo_out[3] = net7;
  assign uo_out[4] = net8;
  assign uo_out[5] = net9;
  assign uo_out[6] = net10;
  assign uo_out[7] = net11;
  assign uio_out[0] = 0;
  assign uio_oe[0] = 0;
  assign uio_out[1] = 0;
  assign uio_oe[1] = 0;
  assign uio_out[2] = 0;
  assign uio_oe[2] = 0;
  assign uio_out[3] = 0;
  assign uio_oe[3] = 0;
  assign uio_out[4] = 0;
  assign uio_oe[4] = 0;
  assign uio_out[5] = 0;
  assign uio_oe[5] = 0;
  assign uio_out[6] = 0;
  assign uio_oe[6] = 0;
  assign uio_out[7] = 0;
  assign uio_oe[7] = 0;

  mux_cell mux1 (
    .a (net17),
    .b (net2),
    .sel (net3),
    .out (net18)
  );
  dff_cell flipflop2 (
    .d (net19),
    .clk (net1),
    .q (net20),
    .notq (net21)
  );
  dff_cell flipflop3 (
    .d (net20),
    .clk (net1),
    .q (net22),
    .notq (net23)
  );
  dff_cell flipflop4 (
    .d (net22),
    .clk (net1),
    .q (net24),
    .notq (net25)
  );
  dff_cell flipflop5 (
    .d (net24),
    .clk (net1),
    .q (net26),
    .notq (net27)
  );
  dff_cell flipflop6 (
    .d (net26),
    .clk (net1),
    .q (net28),
    .notq (net29)
  );
  dff_cell flipflop7 (
    .d (net28),
    .clk (net1),
    .q (net30),
    .notq (net31)
  );
  dff_cell flipflop8 (
    .d (net30),
    .clk (net1),
    .q (net32),
    .notq (net33)
  );
  dff_cell flipflop9 (
    .d (net32),
    .clk (net1),
    .q (net34),
    .notq (net35)
  );
  dff_cell flipflop10 (
    .d (net34),
    .clk (net1),
    .q (net36),
    .notq (net37)
  );
  dff_cell flipflop11 (
    .d (net36),
    .clk (net1),
    .q (net38),
    .notq (net39)
  );
  dff_cell flipflop12 (
    .d (net38),
    .clk (net1),
    .q (net40),
    .notq (net41)
  );
  dff_cell flipflop13 (
    .d (net40),
    .clk (net1),
    .q (net42),
    .notq (net43)
  );
  dff_cell flipflop14 (
    .d (net42),
    .clk (net1),
    .q (net44),
    .notq (net45)
  );
  dff_cell flipflop15 (
    .d (net44),
    .clk (net1),
    .q (net46),
    .notq (net47)
  );
  dff_cell flipflop16 (
    .d (net46),
    .clk (net1),
    .q (net48),
    .notq (net49)
  );
  dff_cell flipflop1 (
    .d (net4),
    .clk (net1),
    .q (net19),
    .notq (net50)
  );
  or_cell gate1 (
    .a (net51),
    .b (net52),
    .out (net17)
  );
  and_cell gate2 (
    .a (net53),
    .b (net54),
    .out (net55)
  );
  and_cell gate4 (
    .a (net21),
    .b (net50),
    .out (net54)
  );
  and_cell gate5 (
    .a (net25),
    .b (net23),
    .out (net53)
  );
  and_cell gate6 (
    .a (net29),
    .b (net27),
    .out (net56)
  );
  and_cell gate9 (
    .a (net33),
    .b (net31),
    .out (net57)
  );
  and_cell gate10 (
    .a (net37),
    .b (net35),
    .out (net58)
  );
  and_cell gate11 (
    .a (net41),
    .b (net39),
    .out (net59)
  );
  and_cell gate12 (
    .a (net45),
    .b (net43),
    .out (net60)
  );
  and_cell gate13 (
    .a (net49),
    .b (net47),
    .out (net61)
  );
  and_cell gate14 (
    .a (net57),
    .b (net56),
    .out (net62)
  );
  and_cell gate15 (
    .a (net59),
    .b (net58),
    .out (net63)
  );
  and_cell gate16 (
    .a (net61),
    .b (net60),
    .out (net64)
  );
  and_cell gate17 (
    .a (net62),
    .b (net55),
    .out (net65)
  );
  and_cell gate19 (
    .a (net64),
    .b (net63),
    .out (net66)
  );
  and_cell gate20 (
    .a (net66),
    .b (net65),
    .out (net67)
  );
  dff_cell flipflop17 (
    .d (net48),
    .clk (net1),
    .q (net68),
    .notq (net69)
  );
  dff_cell flipflop18 (
    .d (net68),
    .clk (net1),
    .q (net70),
    .notq (net71)
  );
  dff_cell flipflop19 (
    .d (net70),
    .clk (net1),
    .q (net72),
    .notq (net73)
  );
  dff_cell flipflop20 (
    .d (net72),
    .clk (net1),
    .q (net74),
    .notq (net75)
  );
  dff_cell flipflop21 (
    .d (net74),
    .clk (net1),
    .q (net76),
    .notq (net77)
  );
  dff_cell flipflop22 (
    .d (net76),
    .clk (net1),
    .q (net78),
    .notq (net79)
  );
  dff_cell flipflop23 (
    .d (net78),
    .clk (net1),
    .q (net80),
    .notq (net81)
  );
  dff_cell flipflop24 (
    .d (net80),
    .clk (net1),
    .q (net82),
    .notq (net83)
  );
  dff_cell flipflop25 (
    .d (net82),
    .clk (net1),
    .q (net84),
    .notq (net85)
  );
  dff_cell flipflop26 (
    .d (net84),
    .clk (net1),
    .q (net86),
    .notq (net87)
  );
  dff_cell flipflop27 (
    .d (net86),
    .clk (net1),
    .q (net88),
    .notq (net89)
  );
  dff_cell flipflop28 (
    .d (net88),
    .clk (net1),
    .q (net90),
    .notq (net91)
  );
  dff_cell flipflop29 (
    .d (net90),
    .clk (net1),
    .q (net92),
    .notq (net93)
  );
  dff_cell flipflop30 (
    .d (net92),
    .clk (net1),
    .q (net94),
    .notq (net95)
  );
  dff_cell flipflop31 (
    .d (net94),
    .clk (net1),
    .q (net96),
    .notq (net97)
  );
  dff_cell flipflop32 (
    .d (net96),
    .clk (net1),
    .q (net98),
    .notq (net99)
  );
  and_cell gate23 (
    .a (net100),
    .b (net101),
    .out (net102)
  );
  and_cell gate24 (
    .a (net71),
    .b (net69),
    .out (net101)
  );
  and_cell gate25 (
    .a (net75),
    .b (net73),
    .out (net100)
  );
  and_cell gate26 (
    .a (net79),
    .b (net77),
    .out (net103)
  );
  and_cell gate32 (
    .a (net81),
    .b (net103),
    .out (net104)
  );
  and_cell gate35 (
    .a (net104),
    .b (net102),
    .out (net105)
  );
  and_cell gate37 (
    .a (net106),
    .b (net105),
    .out (net107)
  );
  and_cell and1 (
    .a (net107),
    .b (net67),
    .out (net108)
  );
  dff_cell flipflop33 (
    .d (net98),
    .clk (net1),
    .q (net109),
    .notq (net110)
  );
  dff_cell flipflop34 (
    .d (net109),
    .clk (net1),
    .q (net111),
    .notq (net112)
  );
  dff_cell flipflop35 (
    .d (net111),
    .clk (net1),
    .q (net113),
    .notq (net114)
  );
  dff_cell flipflop36 (
    .d (net113),
    .clk (net1),
    .q (net115),
    .notq (net116)
  );
  dff_cell flipflop37 (
    .d (net115),
    .clk (net1),
    .q (net117),
    .notq (net118)
  );
  dff_cell flipflop38 (
    .d (net117),
    .clk (net1),
    .q (net119),
    .notq (net120)
  );
  dff_cell flipflop39 (
    .d (net119),
    .clk (net1),
    .q (net121),
    .notq (net122)
  );
  dff_cell flipflop40 (
    .d (net121),
    .clk (net1),
    .q (net123),
    .notq (net124)
  );
  dff_cell flipflop41 (
    .d (net123),
    .clk (net1),
    .q (net125),
    .notq (net126)
  );
  dff_cell flipflop42 (
    .d (net125),
    .clk (net1),
    .q (net127),
    .notq (net128)
  );
  dff_cell flipflop43 (
    .d (net127),
    .clk (net1),
    .q (net129),
    .notq (net130)
  );
  dff_cell flipflop44 (
    .d (net129),
    .clk (net1),
    .q (net131),
    .notq (net132)
  );
  dff_cell flipflop45 (
    .d (net131),
    .clk (net1),
    .q (net133),
    .notq (net134)
  );
  dff_cell flipflop46 (
    .d (net133),
    .clk (net1),
    .q (net135),
    .notq (net136)
  );
  and_cell gate3 (
    .a (net137),
    .b (net138),
    .out (net139)
  );
  and_cell gate7 (
    .a (net85),
    .b (net83),
    .out (net138)
  );
  and_cell gate8 (
    .a (net89),
    .b (net87),
    .out (net137)
  );
  and_cell gate18 (
    .a (net93),
    .b (net91),
    .out (net140)
  );
  and_cell gate21 (
    .a (net97),
    .b (net95),
    .out (net141)
  );
  and_cell gate22 (
    .a (net110),
    .b (net99),
    .out (net142)
  );
  and_cell gate27 (
    .a (net114),
    .b (net112),
    .out (net143)
  );
  and_cell gate28 (
    .a (net118),
    .b (net116),
    .out (net144)
  );
  and_cell gate29 (
    .a (net122),
    .b (net120),
    .out (net145)
  );
  and_cell gate30 (
    .a (net141),
    .b (net140),
    .out (net146)
  );
  and_cell gate31 (
    .a (net143),
    .b (net142),
    .out (net147)
  );
  and_cell gate33 (
    .a (net145),
    .b (net144),
    .out (net148)
  );
  and_cell gate34 (
    .a (net146),
    .b (net139),
    .out (net149)
  );
  and_cell gate36 (
    .a (net148),
    .b (net147),
    .out (net150)
  );
  and_cell gate38 (
    .a (net150),
    .b (net149),
    .out (net151)
  );
  and_cell gate39 (
    .a (net152),
    .b (net153),
    .out (net154)
  );
  and_cell gate40 (
    .a (net126),
    .b (net124),
    .out (net153)
  );
  and_cell gate41 (
    .a (net130),
    .b (net128),
    .out (net152)
  );
  and_cell gate42 (
    .a (net134),
    .b (net132),
    .out (net155)
  );
  and_cell gate43 (
    .a (net136),
    .b (net155),
    .out (net156)
  );
  and_cell gate44 (
    .a (net156),
    .b (net154),
    .out (net106)
  );
  and_cell gate45 (
    .a (net157),
    .b (net151),
    .out (net158)
  );
  dff_cell flipflop47 (
    .d (net135),
    .clk (net1),
    .q (net159),
    .notq (net160)
  );
  dff_cell flipflop48 (
    .d (net159),
    .clk (net1),
    .q (net161),
    .notq (net162)
  );
  dff_cell flipflop49 (
    .d (net161),
    .clk (net1),
    .q (net163),
    .notq (net164)
  );
  dff_cell flipflop50 (
    .d (net163),
    .clk (net1),
    .q (net165),
    .notq (net166)
  );
  dff_cell flipflop51 (
    .d (net165),
    .clk (net1),
    .q (net167),
    .notq (net168)
  );
  dff_cell flipflop52 (
    .d (net167),
    .clk (net1),
    .q (net169),
    .notq (net170)
  );
  dff_cell flipflop53 (
    .d (net169),
    .clk (net1),
    .q (net171),
    .notq (net172)
  );
  dff_cell flipflop54 (
    .d (net171),
    .clk (net1),
    .q (net173),
    .notq (net174)
  );
  dff_cell flipflop55 (
    .d (net173),
    .clk (net1),
    .q (net175),
    .notq (net176)
  );
  dff_cell flipflop56 (
    .d (net175),
    .clk (net1),
    .q (net177),
    .notq (net178)
  );
  dff_cell flipflop57 (
    .d (net177),
    .clk (net1),
    .q (net179),
    .notq (net180)
  );
  dff_cell flipflop58 (
    .d (net179),
    .clk (net1),
    .q (net181),
    .notq (net182)
  );
  dff_cell flipflop59 (
    .d (net181),
    .clk (net1),
    .q (net183),
    .notq (net184)
  );
  dff_cell flipflop60 (
    .d (net183),
    .clk (net1),
    .q (net185),
    .notq (net186)
  );
  dff_cell flipflop61 (
    .d (net185),
    .clk (net1),
    .q (net187),
    .notq (net188)
  );
  dff_cell flipflop62 (
    .d (net187),
    .clk (net1),
    .q (net189),
    .notq (net190)
  );
  and_cell gate46 (
    .a (net191),
    .b (net192),
    .out (net193)
  );
  and_cell gate47 (
    .a (net162),
    .b (net160),
    .out (net192)
  );
  and_cell gate48 (
    .a (net166),
    .b (net164),
    .out (net191)
  );
  and_cell gate49 (
    .a (net170),
    .b (net168),
    .out (net194)
  );
  and_cell gate50 (
    .a (net174),
    .b (net172),
    .out (net195)
  );
  and_cell gate51 (
    .a (net178),
    .b (net176),
    .out (net196)
  );
  and_cell gate52 (
    .a (net182),
    .b (net180),
    .out (net197)
  );
  and_cell gate53 (
    .a (net186),
    .b (net184),
    .out (net198)
  );
  and_cell gate54 (
    .a (net190),
    .b (net188),
    .out (net199)
  );
  and_cell gate55 (
    .a (net195),
    .b (net194),
    .out (net200)
  );
  and_cell gate56 (
    .a (net197),
    .b (net196),
    .out (net201)
  );
  and_cell gate57 (
    .a (net199),
    .b (net198),
    .out (net202)
  );
  and_cell gate58 (
    .a (net200),
    .b (net193),
    .out (net203)
  );
  and_cell gate59 (
    .a (net202),
    .b (net201),
    .out (net204)
  );
  and_cell gate60 (
    .a (net204),
    .b (net203),
    .out (net157)
  );
  dff_cell flipflop63 (
    .d (net189),
    .clk (net1),
    .q (net205),
    .notq (net206)
  );
  dff_cell flipflop64 (
    .d (net205),
    .clk (net1),
    .q (net207),
    .notq (net208)
  );
  dff_cell flipflop65 (
    .d (net207),
    .clk (net1),
    .q (net5),
    .notq (net209)
  );
  dff_cell flipflop66 (
    .d (net5),
    .clk (net1),
    .q (net210),
    .notq (net211)
  );
  dff_cell flipflop67 (
    .d (net210),
    .clk (net1),
    .q (net212),
    .notq (net213)
  );
  dff_cell flipflop68 (
    .d (net212),
    .clk (net1),
    .q (net214),
    .notq (net215)
  );
  dff_cell flipflop69 (
    .d (net214),
    .clk (net1),
    .q (net216),
    .notq (net217)
  );
  dff_cell flipflop70 (
    .d (net216),
    .clk (net1),
    .q (net218),
    .notq (net219)
  );
  dff_cell flipflop71 (
    .d (net218),
    .clk (net1),
    .q (net220),
    .notq (net221)
  );
  dff_cell flipflop72 (
    .d (net220),
    .clk (net1),
    .q (net222),
    .notq (net223)
  );
  dff_cell flipflop73 (
    .d (net222),
    .clk (net1),
    .q (net224),
    .notq (net225)
  );
  dff_cell flipflop74 (
    .d (net224),
    .clk (net1),
    .q (net226),
    .notq (net227)
  );
  dff_cell flipflop75 (
    .d (net226),
    .clk (net1),
    .q (net228),
    .notq (net229)
  );
  dff_cell flipflop76 (
    .d (net228),
    .clk (net1),
    .q (net230),
    .notq (net231)
  );
  dff_cell flipflop77 (
    .d (net230),
    .clk (net1),
    .q (net232),
    .notq (net233)
  );
  dff_cell flipflop78 (
    .d (net232),
    .clk (net1),
    .q (net234),
    .notq (net235)
  );
  and_cell gate61 (
    .a (net236),
    .b (net237),
    .out (net238)
  );
  and_cell gate62 (
    .a (net208),
    .b (net206),
    .out (net237)
  );
  and_cell gate63 (
    .a (net211),
    .b (net209),
    .out (net236)
  );
  and_cell gate64 (
    .a (net215),
    .b (net213),
    .out (net239)
  );
  and_cell gate65 (
    .a (net217),
    .b (net239),
    .out (net240)
  );
  and_cell gate66 (
    .a (net240),
    .b (net238),
    .out (net241)
  );
  and_cell gate67 (
    .a (net242),
    .b (net241),
    .out (net243)
  );
  and_cell and2 (
    .a (net244),
    .b (net243),
    .out (net245)
  );
  dff_cell flipflop79 (
    .d (net234),
    .clk (net1),
    .q (net246),
    .notq (net247)
  );
  dff_cell flipflop80 (
    .d (net246),
    .clk (net1),
    .q (net248),
    .notq (net249)
  );
  dff_cell flipflop81 (
    .d (net248),
    .clk (net1),
    .q (net250),
    .notq (net251)
  );
  dff_cell flipflop82 (
    .d (net250),
    .clk (net1),
    .q (net252),
    .notq (net253)
  );
  dff_cell flipflop83 (
    .d (net252),
    .clk (net1),
    .q (net254),
    .notq (net255)
  );
  dff_cell flipflop84 (
    .d (net254),
    .clk (net1),
    .q (net256),
    .notq (net257)
  );
  dff_cell flipflop85 (
    .d (net256),
    .clk (net1),
    .q (net258),
    .notq (net259)
  );
  dff_cell flipflop86 (
    .d (net258),
    .clk (net1),
    .q (net260),
    .notq (net261)
  );
  dff_cell flipflop87 (
    .d (net260),
    .clk (net1),
    .q (net262),
    .notq (net263)
  );
  dff_cell flipflop88 (
    .d (net262),
    .clk (net1),
    .q (net264),
    .notq (net265)
  );
  dff_cell flipflop89 (
    .d (net264),
    .clk (net1),
    .q (net266),
    .notq (net267)
  );
  dff_cell flipflop90 (
    .d (net266),
    .clk (net1),
    .q (net268),
    .notq (net269)
  );
  dff_cell flipflop91 (
    .d (net268),
    .clk (net1),
    .q (net270),
    .notq (net271)
  );
  dff_cell flipflop92 (
    .d (net270),
    .clk (net1),
    .q (net6),
    .notq (net272)
  );
  and_cell gate68 (
    .a (net273),
    .b (net274),
    .out (net275)
  );
  and_cell gate69 (
    .a (net221),
    .b (net219),
    .out (net274)
  );
  and_cell gate70 (
    .a (net225),
    .b (net223),
    .out (net273)
  );
  and_cell gate71 (
    .a (net229),
    .b (net227),
    .out (net276)
  );
  and_cell gate72 (
    .a (net233),
    .b (net231),
    .out (net277)
  );
  and_cell gate73 (
    .a (net247),
    .b (net235),
    .out (net278)
  );
  and_cell gate74 (
    .a (net251),
    .b (net249),
    .out (net279)
  );
  and_cell gate75 (
    .a (net255),
    .b (net253),
    .out (net280)
  );
  and_cell gate76 (
    .a (net259),
    .b (net257),
    .out (net281)
  );
  and_cell gate77 (
    .a (net277),
    .b (net276),
    .out (net282)
  );
  and_cell gate78 (
    .a (net279),
    .b (net278),
    .out (net283)
  );
  and_cell gate79 (
    .a (net281),
    .b (net280),
    .out (net284)
  );
  and_cell gate80 (
    .a (net282),
    .b (net275),
    .out (net285)
  );
  and_cell gate81 (
    .a (net284),
    .b (net283),
    .out (net286)
  );
  and_cell gate82 (
    .a (net286),
    .b (net285),
    .out (net244)
  );
  and_cell gate83 (
    .a (net287),
    .b (net288),
    .out (net289)
  );
  and_cell gate84 (
    .a (net263),
    .b (net261),
    .out (net288)
  );
  and_cell gate85 (
    .a (net267),
    .b (net265),
    .out (net287)
  );
  and_cell gate86 (
    .a (net271),
    .b (net269),
    .out (net290)
  );
  and_cell gate87 (
    .a (net272),
    .b (net290),
    .out (net291)
  );
  and_cell gate88 (
    .a (net291),
    .b (net289),
    .out (net242)
  );
  and_cell and3 (
    .a (net245),
    .b (net158),
    .out (net292)
  );
  and_cell and4 (
    .a (net292),
    .b (net108),
    .out (net293)
  );
  dff_cell flipflop93 (
    .d (net294),
    .clk (net1),
    .q (net295),
    .notq (net296)
  );
  dff_cell flipflop94 (
    .d (net295),
    .clk (net1),
    .q (net297),
    .notq (net298)
  );
  dff_cell flipflop95 (
    .d (net297),
    .clk (net1),
    .q (net299),
    .notq (net300)
  );
  dff_cell flipflop96 (
    .d (net299),
    .clk (net1),
    .q (net301),
    .notq (net302)
  );
  dff_cell flipflop97 (
    .d (net301),
    .clk (net1),
    .q (net303),
    .notq (net304)
  );
  dff_cell flipflop98 (
    .d (net303),
    .clk (net1),
    .q (net305),
    .notq (net306)
  );
  dff_cell flipflop99 (
    .d (net305),
    .clk (net1),
    .q (net307),
    .notq (net308)
  );
  dff_cell flipflop100 (
    .d (net307),
    .clk (net1),
    .q (net309),
    .notq (net310)
  );
  dff_cell flipflop101 (
    .d (net309),
    .clk (net1),
    .q (net311),
    .notq (net312)
  );
  and_cell gate89 (
    .a (net313),
    .b (net314),
    .out (net315)
  );
  dff_cell flipflop102 (
    .d (net311),
    .clk (net1),
    .q (net316),
    .notq (net317)
  );
  dff_cell flipflop103 (
    .d (net316),
    .clk (net1),
    .q (net318),
    .notq (net319)
  );
  dff_cell flipflop104 (
    .d (net318),
    .clk (net1),
    .q (net320),
    .notq (net321)
  );
  dff_cell flipflop105 (
    .d (net320),
    .clk (net1),
    .q (net322),
    .notq (net323)
  );
  dff_cell flipflop106 (
    .d (net322),
    .clk (net1),
    .q (net324),
    .notq (net325)
  );
  dff_cell flipflop107 (
    .d (net324),
    .clk (net1),
    .q (net326),
    .notq (net327)
  );
  dff_cell flipflop108 (
    .d (net326),
    .clk (net1),
    .q (net328),
    .notq (net329)
  );
  dff_cell flipflop109 (
    .d (net328),
    .clk (net1),
    .q (net330),
    .notq (net331)
  );
  dff_cell flipflop110 (
    .d (net330),
    .clk (net1),
    .q (net332),
    .notq (net333)
  );
  dff_cell flipflop111 (
    .d (net332),
    .clk (net1),
    .q (net334),
    .notq (net335)
  );
  dff_cell flipflop112 (
    .d (net334),
    .clk (net1),
    .q (net336),
    .notq (net337)
  );
  dff_cell flipflop113 (
    .d (net336),
    .clk (net1),
    .q (net338),
    .notq (net339)
  );
  and_cell gate90 (
    .a (net340),
    .b (net341),
    .out (net342)
  );
  and_cell gate91 (
    .a (net298),
    .b (net296),
    .out (net341)
  );
  and_cell gate92 (
    .a (net302),
    .b (net300),
    .out (net340)
  );
  and_cell gate93 (
    .a (net306),
    .b (net304),
    .out (net343)
  );
  and_cell gate94 (
    .a (net310),
    .b (net308),
    .out (net344)
  );
  and_cell gate95 (
    .a (net317),
    .b (net312),
    .out (net345)
  );
  and_cell gate96 (
    .a (net321),
    .b (net319),
    .out (net346)
  );
  and_cell gate97 (
    .a (net325),
    .b (net323),
    .out (net347)
  );
  and_cell gate98 (
    .a (net329),
    .b (net327),
    .out (net348)
  );
  and_cell gate99 (
    .a (net344),
    .b (net343),
    .out (net349)
  );
  and_cell gate100 (
    .a (net346),
    .b (net345),
    .out (net350)
  );
  and_cell gate101 (
    .a (net348),
    .b (net347),
    .out (net351)
  );
  and_cell gate102 (
    .a (net349),
    .b (net342),
    .out (net352)
  );
  and_cell gate103 (
    .a (net351),
    .b (net350),
    .out (net353)
  );
  and_cell gate104 (
    .a (net353),
    .b (net352),
    .out (net354)
  );
  and_cell gate105 (
    .a (net355),
    .b (net356),
    .out (net357)
  );
  and_cell gate106 (
    .a (net333),
    .b (net331),
    .out (net356)
  );
  and_cell gate107 (
    .a (net337),
    .b (net335),
    .out (net355)
  );
  and_cell gate110 (
    .a (net339),
    .b (net357),
    .out (net314)
  );
  dff_cell flipflop114 (
    .d (net338),
    .clk (net1),
    .q (net358),
    .notq (net359)
  );
  dff_cell flipflop115 (
    .d (net358),
    .clk (net1),
    .q (net360),
    .notq (net361)
  );
  dff_cell flipflop116 (
    .d (net360),
    .clk (net1),
    .q (net362),
    .notq (net363)
  );
  dff_cell flipflop117 (
    .d (net362),
    .clk (net1),
    .q (net364),
    .notq (net365)
  );
  dff_cell flipflop118 (
    .d (net364),
    .clk (net1),
    .q (net366),
    .notq (net367)
  );
  dff_cell flipflop119 (
    .d (net366),
    .clk (net1),
    .q (net368),
    .notq (net369)
  );
  dff_cell flipflop120 (
    .d (net368),
    .clk (net1),
    .q (net370),
    .notq (net371)
  );
  dff_cell flipflop121 (
    .d (net370),
    .clk (net1),
    .q (net372),
    .notq (net373)
  );
  dff_cell flipflop122 (
    .d (net372),
    .clk (net1),
    .q (net374),
    .notq (net375)
  );
  dff_cell flipflop123 (
    .d (net374),
    .clk (net1),
    .q (net376),
    .notq (net377)
  );
  dff_cell flipflop124 (
    .d (net376),
    .clk (net1),
    .q (net378),
    .notq (net379)
  );
  dff_cell flipflop125 (
    .d (net378),
    .clk (net1),
    .q (net380),
    .notq (net381)
  );
  dff_cell flipflop126 (
    .d (net380),
    .clk (net1),
    .q (net382),
    .notq (net383)
  );
  dff_cell flipflop127 (
    .d (net382),
    .clk (net1),
    .q (net384),
    .notq (net385)
  );
  dff_cell flipflop128 (
    .d (net384),
    .clk (net1),
    .q (net386),
    .notq (net387)
  );
  dff_cell flipflop129 (
    .d (net386),
    .clk (net1),
    .q (net388),
    .notq (net389)
  );
  dff_cell flipflop130 (
    .d (net388),
    .clk (net1),
    .q (net390),
    .notq (net391)
  );
  dff_cell flipflop131 (
    .d (net390),
    .clk (net1),
    .q (net392),
    .notq (net393)
  );
  dff_cell flipflop132 (
    .d (net392),
    .clk (net1),
    .q (net394),
    .notq (net395)
  );
  dff_cell flipflop133 (
    .d (net394),
    .clk (net1),
    .q (net396),
    .notq (net397)
  );
  dff_cell flipflop134 (
    .d (net396),
    .clk (net1),
    .q (net398),
    .notq (net399)
  );
  and_cell gate109 (
    .a (net400),
    .b (net401),
    .out (net402)
  );
  and_cell gate111 (
    .a (net361),
    .b (net359),
    .out (net401)
  );
  and_cell gate112 (
    .a (net365),
    .b (net363),
    .out (net400)
  );
  and_cell gate113 (
    .a (net369),
    .b (net367),
    .out (net403)
  );
  and_cell gate114 (
    .a (net373),
    .b (net371),
    .out (net404)
  );
  and_cell gate115 (
    .a (net377),
    .b (net375),
    .out (net405)
  );
  and_cell gate116 (
    .a (net381),
    .b (net379),
    .out (net406)
  );
  and_cell gate117 (
    .a (net385),
    .b (net383),
    .out (net407)
  );
  and_cell gate118 (
    .a (net389),
    .b (net387),
    .out (net408)
  );
  and_cell gate119 (
    .a (net404),
    .b (net403),
    .out (net409)
  );
  and_cell gate120 (
    .a (net406),
    .b (net405),
    .out (net410)
  );
  and_cell gate121 (
    .a (net408),
    .b (net407),
    .out (net411)
  );
  and_cell gate122 (
    .a (net409),
    .b (net402),
    .out (net412)
  );
  and_cell gate123 (
    .a (net411),
    .b (net410),
    .out (net413)
  );
  and_cell gate124 (
    .a (net413),
    .b (net412),
    .out (net414)
  );
  and_cell gate125 (
    .a (net415),
    .b (net416),
    .out (net417)
  );
  and_cell gate126 (
    .a (net393),
    .b (net391),
    .out (net416)
  );
  and_cell gate127 (
    .a (net397),
    .b (net395),
    .out (net415)
  );
  and_cell gate128 (
    .a (net399),
    .b (net417),
    .out (net313)
  );
  dff_cell flipflop135 (
    .d (net398),
    .clk (net1),
    .q (net418),
    .notq (net419)
  );
  dff_cell flipflop136 (
    .d (net418),
    .clk (net1),
    .q (net420),
    .notq (net421)
  );
  dff_cell flipflop137 (
    .d (net420),
    .clk (net1),
    .q (net422),
    .notq (net423)
  );
  dff_cell flipflop138 (
    .d (net422),
    .clk (net1),
    .q (net424),
    .notq (net425)
  );
  dff_cell flipflop139 (
    .d (net424),
    .clk (net1),
    .q (net426),
    .notq (net427)
  );
  dff_cell flipflop140 (
    .d (net426),
    .clk (net1),
    .q (net428),
    .notq (net429)
  );
  dff_cell flipflop141 (
    .d (net428),
    .clk (net1),
    .q (net430),
    .notq (net431)
  );
  dff_cell flipflop142 (
    .d (net430),
    .clk (net1),
    .q (net432),
    .notq (net433)
  );
  dff_cell flipflop143 (
    .d (net432),
    .clk (net1),
    .q (net434),
    .notq (net435)
  );
  and_cell gate108 (
    .a (net436),
    .b (net437),
    .out (net438)
  );
  dff_cell flipflop144 (
    .d (net434),
    .clk (net1),
    .q (net439),
    .notq (net440)
  );
  dff_cell flipflop145 (
    .d (net439),
    .clk (net1),
    .q (net441),
    .notq (net442)
  );
  dff_cell flipflop146 (
    .d (net441),
    .clk (net1),
    .q (net443),
    .notq (net444)
  );
  dff_cell flipflop147 (
    .d (net443),
    .clk (net1),
    .q (net445),
    .notq (net446)
  );
  dff_cell flipflop148 (
    .d (net445),
    .clk (net1),
    .q (net447),
    .notq (net448)
  );
  dff_cell flipflop149 (
    .d (net447),
    .clk (net1),
    .q (net449),
    .notq (net450)
  );
  dff_cell flipflop150 (
    .d (net449),
    .clk (net1),
    .q (net451),
    .notq (net452)
  );
  dff_cell flipflop151 (
    .d (net451),
    .clk (net1),
    .q (net453),
    .notq (net454)
  );
  dff_cell flipflop152 (
    .d (net453),
    .clk (net1),
    .q (net455),
    .notq (net456)
  );
  dff_cell flipflop153 (
    .d (net455),
    .clk (net1),
    .q (net457),
    .notq (net458)
  );
  dff_cell flipflop154 (
    .d (net457),
    .clk (net1),
    .q (net459),
    .notq (net460)
  );
  dff_cell flipflop155 (
    .d (net459),
    .clk (net1),
    .q (net461),
    .notq (net462)
  );
  and_cell gate129 (
    .a (net463),
    .b (net464),
    .out (net465)
  );
  and_cell gate130 (
    .a (net421),
    .b (net419),
    .out (net464)
  );
  and_cell gate131 (
    .a (net425),
    .b (net423),
    .out (net463)
  );
  and_cell gate132 (
    .a (net429),
    .b (net427),
    .out (net466)
  );
  and_cell gate133 (
    .a (net433),
    .b (net431),
    .out (net467)
  );
  and_cell gate134 (
    .a (net440),
    .b (net435),
    .out (net468)
  );
  and_cell gate135 (
    .a (net444),
    .b (net442),
    .out (net469)
  );
  and_cell gate136 (
    .a (net448),
    .b (net446),
    .out (net470)
  );
  and_cell gate137 (
    .a (net452),
    .b (net450),
    .out (net471)
  );
  and_cell gate138 (
    .a (net467),
    .b (net466),
    .out (net472)
  );
  and_cell gate139 (
    .a (net469),
    .b (net468),
    .out (net473)
  );
  and_cell gate140 (
    .a (net471),
    .b (net470),
    .out (net474)
  );
  and_cell gate141 (
    .a (net472),
    .b (net465),
    .out (net475)
  );
  and_cell gate142 (
    .a (net474),
    .b (net473),
    .out (net476)
  );
  and_cell gate143 (
    .a (net476),
    .b (net475),
    .out (net477)
  );
  and_cell gate144 (
    .a (net478),
    .b (net479),
    .out (net480)
  );
  and_cell gate145 (
    .a (net456),
    .b (net454),
    .out (net479)
  );
  and_cell gate146 (
    .a (net460),
    .b (net458),
    .out (net478)
  );
  and_cell gate147 (
    .a (net462),
    .b (net480),
    .out (net437)
  );
  dff_cell flipflop156 (
    .d (net461),
    .clk (net1),
    .q (net481),
    .notq (net482)
  );
  dff_cell flipflop157 (
    .d (net481),
    .clk (net1),
    .q (net483),
    .notq (net484)
  );
  dff_cell flipflop158 (
    .d (net483),
    .clk (net1),
    .q (net485),
    .notq (net486)
  );
  dff_cell flipflop159 (
    .d (net485),
    .clk (net1),
    .q (net487),
    .notq (net488)
  );
  dff_cell flipflop160 (
    .d (net487),
    .clk (net1),
    .q (net489),
    .notq (net490)
  );
  dff_cell flipflop161 (
    .d (net489),
    .clk (net1),
    .q (net7),
    .notq (net491)
  );
  dff_cell flipflop162 (
    .d (net7),
    .clk (net1),
    .q (net492),
    .notq (net493)
  );
  dff_cell flipflop163 (
    .d (net492),
    .clk (net1),
    .q (net494),
    .notq (net495)
  );
  dff_cell flipflop164 (
    .d (net494),
    .clk (net1),
    .q (net496),
    .notq (net497)
  );
  dff_cell flipflop165 (
    .d (net496),
    .clk (net1),
    .q (net498),
    .notq (net499)
  );
  dff_cell flipflop166 (
    .d (net498),
    .clk (net1),
    .q (net500),
    .notq (net501)
  );
  dff_cell flipflop167 (
    .d (net500),
    .clk (net1),
    .q (net502),
    .notq (net503)
  );
  dff_cell flipflop168 (
    .d (net502),
    .clk (net1),
    .q (net504),
    .notq (net505)
  );
  dff_cell flipflop169 (
    .d (net504),
    .clk (net1),
    .q (net506),
    .notq (net507)
  );
  dff_cell flipflop170 (
    .d (net506),
    .clk (net1),
    .q (net508),
    .notq (net509)
  );
  dff_cell flipflop171 (
    .d (net508),
    .clk (net1),
    .q (net510),
    .notq (net511)
  );
  dff_cell flipflop172 (
    .d (net510),
    .clk (net1),
    .q (net512),
    .notq (net513)
  );
  dff_cell flipflop173 (
    .d (net512),
    .clk (net1),
    .q (net514),
    .notq (net515)
  );
  dff_cell flipflop174 (
    .d (net514),
    .clk (net1),
    .q (net516),
    .notq (net517)
  );
  dff_cell flipflop175 (
    .d (net516),
    .clk (net1),
    .q (net518),
    .notq (net519)
  );
  dff_cell flipflop176 (
    .d (net518),
    .clk (net1),
    .q (net8),
    .notq (net520)
  );
  and_cell gate148 (
    .a (net521),
    .b (net522),
    .out (net523)
  );
  and_cell gate149 (
    .a (net484),
    .b (net482),
    .out (net522)
  );
  and_cell gate150 (
    .a (net488),
    .b (net486),
    .out (net521)
  );
  and_cell gate151 (
    .a (net491),
    .b (net490),
    .out (net524)
  );
  and_cell gate152 (
    .a (net495),
    .b (net493),
    .out (net525)
  );
  and_cell gate153 (
    .a (net499),
    .b (net497),
    .out (net526)
  );
  and_cell gate154 (
    .a (net503),
    .b (net501),
    .out (net527)
  );
  and_cell gate155 (
    .a (net507),
    .b (net505),
    .out (net528)
  );
  and_cell gate156 (
    .a (net511),
    .b (net509),
    .out (net529)
  );
  and_cell gate157 (
    .a (net525),
    .b (net524),
    .out (net530)
  );
  and_cell gate158 (
    .a (net527),
    .b (net526),
    .out (net531)
  );
  and_cell gate159 (
    .a (net529),
    .b (net528),
    .out (net532)
  );
  and_cell gate160 (
    .a (net530),
    .b (net523),
    .out (net533)
  );
  and_cell gate161 (
    .a (net532),
    .b (net531),
    .out (net534)
  );
  and_cell gate162 (
    .a (net534),
    .b (net533),
    .out (net535)
  );
  and_cell gate163 (
    .a (net536),
    .b (net537),
    .out (net538)
  );
  and_cell gate164 (
    .a (net515),
    .b (net513),
    .out (net537)
  );
  and_cell gate165 (
    .a (net519),
    .b (net517),
    .out (net536)
  );
  and_cell gate166 (
    .a (net520),
    .b (net538),
    .out (net436)
  );
  and_cell gate167 (
    .a (net315),
    .b (net354),
    .out (net539)
  );
  and_cell gate168 (
    .a (net414),
    .b (net539),
    .out (net540)
  );
  and_cell gate169 (
    .a (net438),
    .b (net477),
    .out (net541)
  );
  and_cell gate170 (
    .a (net535),
    .b (net541),
    .out (net542)
  );
  and_cell gate171 (
    .a (net542),
    .b (net540),
    .out (net543)
  );
  and_cell gate172 (
    .a (net543),
    .b (net293),
    .out (net544)
  );
  dff_cell flipflop0 (
    .d (net18),
    .clk (net1),
    .q (net4),
    .notq (net545)
  );
  and_cell gate173 (
    .a (net544),
    .b (net545),
    .out (net546)
  );
  and_cell and5 (
    .a (net268),
    .b (net270),
    .out (net547)
  );
  xor_cell xor1 (
    .a (net6),
    .b (net5),
    .out (net548)
  );
  xor_cell xor2 (
    .a (net548),
    .b (net547),
    .out (net549)
  );
  xor_cell xor3 (
    .a (net508),
    .b (net549),
    .out (net550)
  );
  mux_cell mux2 (
    .a (net550),
    .b (net6),
    .sel (net3),
    .out (net294)
  );
  and_cell and6 (
    .a (net516),
    .b (net518),
    .out (net551)
  );
  xor_cell xor4 (
    .a (net8),
    .b (net7),
    .out (net552)
  );
  xor_cell xor5 (
    .a (net552),
    .b (net551),
    .out (net553)
  );
  xor_cell xor6 (
    .a (net552),
    .b (net548),
    .out (net554)
  );
  xor_cell xor7 (
    .a (net555),
    .b (net214),
    .out (net52)
  );
  dff_cell flipflop177 (
    .d (net556),
    .clk (net1),
    .q (net557),
    .notq (net558)
  );
  dff_cell flipflop178 (
    .d (net557),
    .clk (net1),
    .q (net559),
    .notq (net560)
  );
  dff_cell flipflop179 (
    .d (net559),
    .clk (net1),
    .q (net561),
    .notq (net562)
  );
  dff_cell flipflop180 (
    .d (net561),
    .clk (net1),
    .q (net563),
    .notq (net564)
  );
  dff_cell flipflop181 (
    .d (net563),
    .clk (net1),
    .q (net565),
    .notq (net566)
  );
  dff_cell flipflop182 (
    .d (net565),
    .clk (net1),
    .q (net567),
    .notq (net568)
  );
  dff_cell flipflop183 (
    .d (net567),
    .clk (net1),
    .q (net569),
    .notq (net570)
  );
  dff_cell flipflop184 (
    .d (net569),
    .clk (net1),
    .q (net571),
    .notq (net572)
  );
  dff_cell flipflop185 (
    .d (net571),
    .clk (net1),
    .q (net573),
    .notq (net574)
  );
  dff_cell flipflop186 (
    .d (net573),
    .clk (net1),
    .q (net575),
    .notq (net576)
  );
  dff_cell flipflop187 (
    .d (net575),
    .clk (net1),
    .q (net577),
    .notq (net578)
  );
  dff_cell flipflop188 (
    .d (net577),
    .clk (net1),
    .q (net579),
    .notq (net580)
  );
  dff_cell flipflop189 (
    .d (net579),
    .clk (net1),
    .q (net581),
    .notq (net582)
  );
  dff_cell flipflop190 (
    .d (net581),
    .clk (net1),
    .q (net583),
    .notq (net584)
  );
  dff_cell flipflop191 (
    .d (net583),
    .clk (net1),
    .q (net585),
    .notq (net586)
  );
  dff_cell flipflop192 (
    .d (net585),
    .clk (net1),
    .q (net587),
    .notq (net588)
  );
  dff_cell flipflop193 (
    .d (net587),
    .clk (net1),
    .q (net589),
    .notq (net590)
  );
  dff_cell flipflop194 (
    .d (net589),
    .clk (net1),
    .q (net591),
    .notq (net592)
  );
  dff_cell flipflop195 (
    .d (net591),
    .clk (net1),
    .q (net593),
    .notq (net594)
  );
  dff_cell flipflop196 (
    .d (net593),
    .clk (net1),
    .q (net595),
    .notq (net596)
  );
  dff_cell flipflop197 (
    .d (net595),
    .clk (net1),
    .q (net597),
    .notq (net598)
  );
  and_cell gate174 (
    .a (net599),
    .b (net600),
    .out (net601)
  );
  and_cell gate175 (
    .a (net560),
    .b (net558),
    .out (net600)
  );
  and_cell gate176 (
    .a (net564),
    .b (net562),
    .out (net599)
  );
  and_cell gate177 (
    .a (net568),
    .b (net566),
    .out (net602)
  );
  and_cell gate178 (
    .a (net572),
    .b (net570),
    .out (net603)
  );
  and_cell gate179 (
    .a (net576),
    .b (net574),
    .out (net604)
  );
  and_cell gate180 (
    .a (net580),
    .b (net578),
    .out (net605)
  );
  and_cell gate181 (
    .a (net584),
    .b (net582),
    .out (net606)
  );
  and_cell gate182 (
    .a (net588),
    .b (net586),
    .out (net607)
  );
  and_cell gate183 (
    .a (net592),
    .b (net590),
    .out (net608)
  );
  and_cell gate184 (
    .a (net596),
    .b (net594),
    .out (net609)
  );
  dff_cell flipflop198 (
    .d (net597),
    .clk (net1),
    .q (net610),
    .notq (net611)
  );
  and_cell gate185 (
    .a (net611),
    .b (net598),
    .out (net612)
  );
  and_cell gate186 (
    .a (net603),
    .b (net602),
    .out (net613)
  );
  and_cell gate187 (
    .a (net605),
    .b (net604),
    .out (net614)
  );
  and_cell gate188 (
    .a (net607),
    .b (net606),
    .out (net615)
  );
  and_cell gate189 (
    .a (net609),
    .b (net608),
    .out (net616)
  );
  and_cell gate190 (
    .a (net613),
    .b (net601),
    .out (net617)
  );
  and_cell gate191 (
    .a (net615),
    .b (net614),
    .out (net618)
  );
  dff_cell flipflop199 (
    .d (net610),
    .clk (net1),
    .q (net619),
    .notq (net620)
  );
  dff_cell flipflop200 (
    .d (net619),
    .clk (net1),
    .q (net621),
    .notq (net622)
  );
  dff_cell flipflop201 (
    .d (net621),
    .clk (net1),
    .q (net623),
    .notq (net624)
  );
  dff_cell flipflop202 (
    .d (net623),
    .clk (net1),
    .q (net625),
    .notq (net626)
  );
  dff_cell flipflop203 (
    .d (net625),
    .clk (net1),
    .q (net627),
    .notq (net628)
  );
  dff_cell flipflop204 (
    .d (net627),
    .clk (net1),
    .q (net629),
    .notq (net630)
  );
  dff_cell flipflop205 (
    .d (net629),
    .clk (net1),
    .q (net631),
    .notq (net632)
  );
  dff_cell flipflop206 (
    .d (net631),
    .clk (net1),
    .q (net633),
    .notq (net634)
  );
  dff_cell flipflop207 (
    .d (net633),
    .clk (net1),
    .q (net635),
    .notq (net636)
  );
  dff_cell flipflop208 (
    .d (net635),
    .clk (net1),
    .q (net637),
    .notq (net638)
  );
  dff_cell flipflop209 (
    .d (net637),
    .clk (net1),
    .q (net639),
    .notq (net640)
  );
  dff_cell flipflop210 (
    .d (net639),
    .clk (net1),
    .q (net641),
    .notq (net642)
  );
  dff_cell flipflop211 (
    .d (net641),
    .clk (net1),
    .q (net643),
    .notq (net644)
  );
  dff_cell flipflop212 (
    .d (net643),
    .clk (net1),
    .q (net645),
    .notq (net646)
  );
  dff_cell flipflop213 (
    .d (net645),
    .clk (net1),
    .q (net647),
    .notq (net648)
  );
  dff_cell flipflop214 (
    .d (net647),
    .clk (net1),
    .q (net649),
    .notq (net650)
  );
  dff_cell flipflop215 (
    .d (net649),
    .clk (net1),
    .q (net651),
    .notq (net652)
  );
  dff_cell flipflop216 (
    .d (net651),
    .clk (net1),
    .q (net653),
    .notq (net654)
  );
  dff_cell flipflop217 (
    .d (net653),
    .clk (net1),
    .q (net655),
    .notq (net656)
  );
  dff_cell flipflop218 (
    .d (net655),
    .clk (net1),
    .q (net657),
    .notq (net658)
  );
  dff_cell flipflop219 (
    .d (net657),
    .clk (net1),
    .q (net659),
    .notq (net660)
  );
  and_cell gate192 (
    .a (net661),
    .b (net662),
    .out (net663)
  );
  and_cell gate193 (
    .a (net622),
    .b (net620),
    .out (net662)
  );
  and_cell gate194 (
    .a (net626),
    .b (net624),
    .out (net661)
  );
  and_cell gate195 (
    .a (net630),
    .b (net628),
    .out (net664)
  );
  and_cell gate196 (
    .a (net634),
    .b (net632),
    .out (net665)
  );
  and_cell gate197 (
    .a (net638),
    .b (net636),
    .out (net666)
  );
  and_cell gate198 (
    .a (net642),
    .b (net640),
    .out (net667)
  );
  and_cell gate199 (
    .a (net646),
    .b (net644),
    .out (net668)
  );
  and_cell gate200 (
    .a (net650),
    .b (net648),
    .out (net669)
  );
  and_cell gate201 (
    .a (net654),
    .b (net652),
    .out (net670)
  );
  and_cell gate202 (
    .a (net658),
    .b (net656),
    .out (net671)
  );
  dff_cell flipflop220 (
    .d (net659),
    .clk (net1),
    .q (net672),
    .notq (net673)
  );
  and_cell gate203 (
    .a (net673),
    .b (net660),
    .out (net674)
  );
  and_cell gate204 (
    .a (net665),
    .b (net664),
    .out (net675)
  );
  and_cell gate205 (
    .a (net667),
    .b (net666),
    .out (net676)
  );
  and_cell gate206 (
    .a (net669),
    .b (net668),
    .out (net677)
  );
  and_cell gate207 (
    .a (net671),
    .b (net670),
    .out (net678)
  );
  and_cell gate208 (
    .a (net675),
    .b (net663),
    .out (net679)
  );
  and_cell gate209 (
    .a (net677),
    .b (net676),
    .out (net680)
  );
  dff_cell flipflop221 (
    .d (net672),
    .clk (net1),
    .q (net681),
    .notq (net682)
  );
  dff_cell flipflop222 (
    .d (net681),
    .clk (net1),
    .q (net683),
    .notq (net684)
  );
  dff_cell flipflop223 (
    .d (net683),
    .clk (net1),
    .q (net685),
    .notq (net686)
  );
  dff_cell flipflop224 (
    .d (net685),
    .clk (net1),
    .q (net687),
    .notq (net688)
  );
  dff_cell flipflop225 (
    .d (net687),
    .clk (net1),
    .q (net689),
    .notq (net690)
  );
  dff_cell flipflop226 (
    .d (net689),
    .clk (net1),
    .q (net691),
    .notq (net692)
  );
  dff_cell flipflop227 (
    .d (net691),
    .clk (net1),
    .q (net693),
    .notq (net694)
  );
  dff_cell flipflop228 (
    .d (net693),
    .clk (net1),
    .q (net695),
    .notq (net696)
  );
  dff_cell flipflop229 (
    .d (net695),
    .clk (net1),
    .q (net697),
    .notq (net698)
  );
  dff_cell flipflop230 (
    .d (net697),
    .clk (net1),
    .q (net699),
    .notq (net700)
  );
  dff_cell flipflop231 (
    .d (net699),
    .clk (net1),
    .q (net701),
    .notq (net702)
  );
  dff_cell flipflop232 (
    .d (net701),
    .clk (net1),
    .q (net703),
    .notq (net704)
  );
  dff_cell flipflop233 (
    .d (net703),
    .clk (net1),
    .q (net705),
    .notq (net706)
  );
  dff_cell flipflop234 (
    .d (net705),
    .clk (net1),
    .q (net707),
    .notq (net708)
  );
  dff_cell flipflop235 (
    .d (net707),
    .clk (net1),
    .q (net709),
    .notq (net710)
  );
  dff_cell flipflop236 (
    .d (net709),
    .clk (net1),
    .q (net711),
    .notq (net712)
  );
  dff_cell flipflop237 (
    .d (net711),
    .clk (net1),
    .q (net713),
    .notq (net714)
  );
  dff_cell flipflop238 (
    .d (net713),
    .clk (net1),
    .q (net715),
    .notq (net716)
  );
  dff_cell flipflop239 (
    .d (net715),
    .clk (net1),
    .q (net717),
    .notq (net718)
  );
  dff_cell flipflop240 (
    .d (net717),
    .clk (net1),
    .q (net719),
    .notq (net720)
  );
  dff_cell flipflop241 (
    .d (net719),
    .clk (net1),
    .q (net721),
    .notq (net722)
  );
  and_cell gate210 (
    .a (net723),
    .b (net724),
    .out (net725)
  );
  and_cell gate211 (
    .a (net684),
    .b (net682),
    .out (net724)
  );
  and_cell gate212 (
    .a (net688),
    .b (net686),
    .out (net723)
  );
  and_cell gate213 (
    .a (net692),
    .b (net690),
    .out (net726)
  );
  and_cell gate214 (
    .a (net696),
    .b (net694),
    .out (net727)
  );
  and_cell gate215 (
    .a (net700),
    .b (net698),
    .out (net728)
  );
  and_cell gate216 (
    .a (net704),
    .b (net702),
    .out (net729)
  );
  and_cell gate217 (
    .a (net708),
    .b (net706),
    .out (net730)
  );
  and_cell gate218 (
    .a (net712),
    .b (net710),
    .out (net731)
  );
  and_cell gate219 (
    .a (net716),
    .b (net714),
    .out (net732)
  );
  and_cell gate220 (
    .a (net720),
    .b (net718),
    .out (net733)
  );
  dff_cell flipflop242 (
    .d (net721),
    .clk (net1),
    .q (net9),
    .notq (net734)
  );
  and_cell gate221 (
    .a (net734),
    .b (net722),
    .out (net735)
  );
  and_cell gate222 (
    .a (net727),
    .b (net726),
    .out (net736)
  );
  and_cell gate223 (
    .a (net729),
    .b (net728),
    .out (net737)
  );
  and_cell gate224 (
    .a (net731),
    .b (net730),
    .out (net738)
  );
  and_cell gate225 (
    .a (net733),
    .b (net732),
    .out (net739)
  );
  and_cell gate226 (
    .a (net736),
    .b (net725),
    .out (net740)
  );
  and_cell gate227 (
    .a (net738),
    .b (net737),
    .out (net741)
  );
  dff_cell flipflop243 (
    .d (net9),
    .clk (net1),
    .q (net742),
    .notq (net743)
  );
  dff_cell flipflop244 (
    .d (net742),
    .clk (net1),
    .q (net744),
    .notq (net745)
  );
  dff_cell flipflop245 (
    .d (net744),
    .clk (net1),
    .q (net746),
    .notq (net747)
  );
  dff_cell flipflop246 (
    .d (net746),
    .clk (net1),
    .q (net748),
    .notq (net749)
  );
  dff_cell flipflop247 (
    .d (net748),
    .clk (net1),
    .q (net750),
    .notq (net751)
  );
  dff_cell flipflop248 (
    .d (net750),
    .clk (net1),
    .q (net752),
    .notq (net753)
  );
  dff_cell flipflop249 (
    .d (net752),
    .clk (net1),
    .q (net754),
    .notq (net755)
  );
  dff_cell flipflop250 (
    .d (net754),
    .clk (net1),
    .q (net756),
    .notq (net757)
  );
  dff_cell flipflop251 (
    .d (net756),
    .clk (net1),
    .q (net758),
    .notq (net759)
  );
  dff_cell flipflop252 (
    .d (net758),
    .clk (net1),
    .q (net760),
    .notq (net761)
  );
  dff_cell flipflop253 (
    .d (net760),
    .clk (net1),
    .q (net762),
    .notq (net763)
  );
  dff_cell flipflop254 (
    .d (net762),
    .clk (net1),
    .q (net764),
    .notq (net765)
  );
  dff_cell flipflop255 (
    .d (net764),
    .clk (net1),
    .q (net766),
    .notq (net767)
  );
  dff_cell flipflop256 (
    .d (net766),
    .clk (net1),
    .q (net768),
    .notq (net769)
  );
  dff_cell flipflop257 (
    .d (net768),
    .clk (net1),
    .q (net770),
    .notq (net771)
  );
  dff_cell flipflop258 (
    .d (net770),
    .clk (net1),
    .q (net772),
    .notq (net773)
  );
  dff_cell flipflop259 (
    .d (net772),
    .clk (net1),
    .q (net774),
    .notq (net775)
  );
  dff_cell flipflop260 (
    .d (net774),
    .clk (net1),
    .q (net776),
    .notq (net777)
  );
  dff_cell flipflop261 (
    .d (net776),
    .clk (net1),
    .q (net778),
    .notq (net779)
  );
  dff_cell flipflop262 (
    .d (net778),
    .clk (net1),
    .q (net780),
    .notq (net781)
  );
  dff_cell flipflop263 (
    .d (net780),
    .clk (net1),
    .q (net782),
    .notq (net783)
  );
  and_cell gate228 (
    .a (net784),
    .b (net785),
    .out (net786)
  );
  and_cell gate229 (
    .a (net745),
    .b (net743),
    .out (net785)
  );
  and_cell gate230 (
    .a (net749),
    .b (net747),
    .out (net784)
  );
  and_cell gate231 (
    .a (net753),
    .b (net751),
    .out (net787)
  );
  and_cell gate232 (
    .a (net757),
    .b (net755),
    .out (net788)
  );
  and_cell gate233 (
    .a (net761),
    .b (net759),
    .out (net789)
  );
  and_cell gate234 (
    .a (net765),
    .b (net763),
    .out (net790)
  );
  and_cell gate235 (
    .a (net769),
    .b (net767),
    .out (net791)
  );
  and_cell gate236 (
    .a (net773),
    .b (net771),
    .out (net792)
  );
  and_cell gate237 (
    .a (net777),
    .b (net775),
    .out (net793)
  );
  and_cell gate238 (
    .a (net781),
    .b (net779),
    .out (net794)
  );
  dff_cell flipflop264 (
    .d (net782),
    .clk (net1),
    .q (net795),
    .notq (net796)
  );
  and_cell gate239 (
    .a (net796),
    .b (net783),
    .out (net797)
  );
  and_cell gate240 (
    .a (net788),
    .b (net787),
    .out (net798)
  );
  and_cell gate241 (
    .a (net790),
    .b (net789),
    .out (net799)
  );
  and_cell gate242 (
    .a (net792),
    .b (net791),
    .out (net800)
  );
  and_cell gate243 (
    .a (net794),
    .b (net793),
    .out (net801)
  );
  and_cell gate244 (
    .a (net798),
    .b (net786),
    .out (net802)
  );
  and_cell gate245 (
    .a (net800),
    .b (net799),
    .out (net803)
  );
  dff_cell flipflop265 (
    .d (net795),
    .clk (net1),
    .q (net804),
    .notq (net805)
  );
  dff_cell flipflop266 (
    .d (net804),
    .clk (net1),
    .q (net806),
    .notq (net807)
  );
  dff_cell flipflop267 (
    .d (net806),
    .clk (net1),
    .q (net808),
    .notq (net809)
  );
  dff_cell flipflop268 (
    .d (net808),
    .clk (net1),
    .q (net810),
    .notq (net811)
  );
  dff_cell flipflop269 (
    .d (net810),
    .clk (net1),
    .q (net812),
    .notq (net813)
  );
  dff_cell flipflop270 (
    .d (net812),
    .clk (net1),
    .q (net814),
    .notq (net815)
  );
  dff_cell flipflop271 (
    .d (net814),
    .clk (net1),
    .q (net816),
    .notq (net817)
  );
  dff_cell flipflop272 (
    .d (net816),
    .clk (net1),
    .q (net818),
    .notq (net819)
  );
  dff_cell flipflop273 (
    .d (net818),
    .clk (net1),
    .q (net820),
    .notq (net821)
  );
  dff_cell flipflop274 (
    .d (net820),
    .clk (net1),
    .q (net822),
    .notq (net823)
  );
  dff_cell flipflop275 (
    .d (net822),
    .clk (net1),
    .q (net824),
    .notq (net825)
  );
  dff_cell flipflop276 (
    .d (net824),
    .clk (net1),
    .q (net826),
    .notq (net827)
  );
  dff_cell flipflop277 (
    .d (net826),
    .clk (net1),
    .q (net828),
    .notq (net829)
  );
  dff_cell flipflop278 (
    .d (net828),
    .clk (net1),
    .q (net830),
    .notq (net831)
  );
  dff_cell flipflop279 (
    .d (net830),
    .clk (net1),
    .q (net832),
    .notq (net833)
  );
  dff_cell flipflop280 (
    .d (net832),
    .clk (net1),
    .q (net834),
    .notq (net835)
  );
  dff_cell flipflop281 (
    .d (net834),
    .clk (net1),
    .q (net836),
    .notq (net837)
  );
  dff_cell flipflop282 (
    .d (net836),
    .clk (net1),
    .q (net838),
    .notq (net839)
  );
  dff_cell flipflop283 (
    .d (net838),
    .clk (net1),
    .q (net840),
    .notq (net841)
  );
  dff_cell flipflop284 (
    .d (net840),
    .clk (net1),
    .q (net842),
    .notq (net843)
  );
  dff_cell flipflop285 (
    .d (net842),
    .clk (net1),
    .q (net844),
    .notq (net845)
  );
  and_cell gate246 (
    .a (net846),
    .b (net847),
    .out (net848)
  );
  and_cell gate247 (
    .a (net807),
    .b (net805),
    .out (net847)
  );
  and_cell gate248 (
    .a (net811),
    .b (net809),
    .out (net846)
  );
  and_cell gate249 (
    .a (net815),
    .b (net813),
    .out (net849)
  );
  and_cell gate250 (
    .a (net819),
    .b (net817),
    .out (net850)
  );
  and_cell gate251 (
    .a (net823),
    .b (net821),
    .out (net851)
  );
  and_cell gate252 (
    .a (net827),
    .b (net825),
    .out (net852)
  );
  and_cell gate253 (
    .a (net831),
    .b (net829),
    .out (net853)
  );
  and_cell gate254 (
    .a (net835),
    .b (net833),
    .out (net854)
  );
  and_cell gate255 (
    .a (net839),
    .b (net837),
    .out (net855)
  );
  and_cell gate256 (
    .a (net843),
    .b (net841),
    .out (net856)
  );
  dff_cell flipflop286 (
    .d (net844),
    .clk (net1),
    .q (net857),
    .notq (net858)
  );
  and_cell gate257 (
    .a (net858),
    .b (net845),
    .out (net859)
  );
  and_cell gate258 (
    .a (net850),
    .b (net849),
    .out (net860)
  );
  and_cell gate259 (
    .a (net852),
    .b (net851),
    .out (net861)
  );
  and_cell gate260 (
    .a (net854),
    .b (net853),
    .out (net862)
  );
  and_cell gate261 (
    .a (net856),
    .b (net855),
    .out (net863)
  );
  and_cell gate262 (
    .a (net860),
    .b (net848),
    .out (net864)
  );
  and_cell gate263 (
    .a (net862),
    .b (net861),
    .out (net865)
  );
  dff_cell flipflop287 (
    .d (net857),
    .clk (net1),
    .q (net10),
    .notq (net866)
  );
  and_cell gate264 (
    .a (net612),
    .b (net616),
    .out (net867)
  );
  and_cell gate265 (
    .a (net674),
    .b (net678),
    .out (net868)
  );
  and_cell gate266 (
    .a (net735),
    .b (net739),
    .out (net869)
  );
  and_cell gate267 (
    .a (net797),
    .b (net801),
    .out (net870)
  );
  and_cell gate268 (
    .a (net859),
    .b (net863),
    .out (net871)
  );
  and_cell gate269 (
    .a (net866),
    .b (net871),
    .out (net872)
  );
  and_cell gate270 (
    .a (net618),
    .b (net617),
    .out (net873)
  );
  and_cell gate271 (
    .a (net679),
    .b (net867),
    .out (net874)
  );
  and_cell gate272 (
    .a (net868),
    .b (net680),
    .out (net875)
  );
  and_cell gate273 (
    .a (net741),
    .b (net740),
    .out (net876)
  );
  and_cell gate274 (
    .a (net802),
    .b (net869),
    .out (net877)
  );
  and_cell gate275 (
    .a (net870),
    .b (net803),
    .out (net878)
  );
  and_cell gate276 (
    .a (net865),
    .b (net864),
    .out (net879)
  );
  and_cell gate277 (
    .a (net872),
    .b (net879),
    .out (net880)
  );
  and_cell gate278 (
    .a (net880),
    .b (net878),
    .out (net881)
  );
  and_cell gate279 (
    .a (net877),
    .b (net876),
    .out (net882)
  );
  and_cell gate280 (
    .a (net874),
    .b (net873),
    .out (net883)
  );
  and_cell gate281 (
    .a (net882),
    .b (net875),
    .out (net884)
  );
  and_cell gate282 (
    .a (net884),
    .b (net883),
    .out (net885)
  );
  and_cell gate283 (
    .a (net881),
    .b (net885),
    .out (net886)
  );
  and_cell and7 (
    .a (net546),
    .b (net886),
    .out (net51)
  );
  xor_cell xor8 (
    .a (net782),
    .b (net553),
    .out (net887)
  );
  and_cell and8 (
    .a (net857),
    .b (net844),
    .out (net888)
  );
  xor_cell xor9 (
    .a (net10),
    .b (net9),
    .out (net889)
  );
  xor_cell xor10 (
    .a (net889),
    .b (net888),
    .out (net555)
  );
  xor_cell xor11 (
    .a (net554),
    .b (net889),
    .out (net11)
  );
  mux_cell mux3 (
    .a (net887),
    .b (net8),
    .sel (net3),
    .out (net556)
  );
endmodule
