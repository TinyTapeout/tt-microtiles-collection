/* Automatically generated from https://wokwi.com/projects/395263962779770881 */

`default_nettype none

module tt_um_wokwi_395263962779770881(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = ui_in[1];
  wire net3 = ui_in[2];
  wire net4;
  wire net5;
  wire net6;
  wire net7;
  wire net8;
  wire net9;
  wire net10;
  wire net11;
  wire net12 = 1'b0;
  wire net13 = 1'b1;
  wire net14 = 1'b1;
  wire net15 = 1'b0;
  wire net16 = 1'b1;
  wire net17;
  wire net18;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291;
  wire net292;
  wire net293;
  wire net294;
  wire net295;
  wire net296;
  wire net297;
  wire net298;
  wire net299;
  wire net300;
  wire net301;
  wire net302;
  wire net303;
  wire net304;
  wire net305;
  wire net306;
  wire net307;
  wire net308;
  wire net309;
  wire net310;
  wire net311;
  wire net312;
  wire net313;
  wire net314;
  wire net315;
  wire net316;
  wire net317;
  wire net318;
  wire net319;
  wire net320;
  wire net321;
  wire net322;
  wire net323;
  wire net324;
  wire net325;
  wire net326;
  wire net327;
  wire net328;
  wire net329;
  wire net330;
  wire net331;
  wire net332;
  wire net333;
  wire net334;
  wire net335;
  wire net336;
  wire net337;
  wire net338;
  wire net339;
  wire net340;
  wire net341;
  wire net342;
  wire net343;
  wire net344;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349;
  wire net350;
  wire net351;
  wire net352;
  wire net353;
  wire net354;
  wire net355;
  wire net356;
  wire net357;
  wire net358;
  wire net359;
  wire net360;
  wire net361;
  wire net362;
  wire net363;
  wire net364;
  wire net365;
  wire net366;
  wire net367;
  wire net368;
  wire net369;
  wire net370;
  wire net371;
  wire net372;
  wire net373;
  wire net374;
  wire net375;
  wire net376;
  wire net377;
  wire net378;
  wire net379;
  wire net380;
  wire net381;
  wire net382;
  wire net383;
  wire net384;
  wire net385;
  wire net386;
  wire net387;
  wire net388;
  wire net389;
  wire net390;
  wire net391;
  wire net392;
  wire net393;
  wire net394;
  wire net395;
  wire net396;
  wire net397;
  wire net398;
  wire net399;
  wire net400;
  wire net401;
  wire net402;
  wire net403;
  wire net404;
  wire net405;
  wire net406;
  wire net407;
  wire net408;
  wire net409;
  wire net410;
  wire net411;
  wire net412;
  wire net413;
  wire net414;
  wire net415;
  wire net416;
  wire net417;
  wire net418;
  wire net419;
  wire net420;
  wire net421;
  wire net422;
  wire net423;
  wire net424;
  wire net425;
  wire net426;
  wire net427;
  wire net428;
  wire net429;
  wire net430;
  wire net431;
  wire net432;
  wire net433;
  wire net434;
  wire net435;
  wire net436;
  wire net437;
  wire net438;
  wire net439;
  wire net440;
  wire net441;
  wire net442;
  wire net443;
  wire net444;
  wire net445;
  wire net446;
  wire net447;
  wire net448;
  wire net449;
  wire net450;
  wire net451;
  wire net452;
  wire net453;
  wire net454;
  wire net455;
  wire net456;
  wire net457;
  wire net458;
  wire net459;
  wire net460;
  wire net461;
  wire net462;
  wire net463;
  wire net464;
  wire net465;
  wire net466;
  wire net467;
  wire net468;
  wire net469;
  wire net470;
  wire net471;
  wire net472;
  wire net473;
  wire net474;
  wire net475;
  wire net476;
  wire net477;
  wire net478;
  wire net479;
  wire net480;
  wire net481;
  wire net482;
  wire net483;
  wire net484;
  wire net485;
  wire net486;
  wire net487;
  wire net488;
  wire net489;
  wire net490;
  wire net491;
  wire net492;
  wire net493;
  wire net494;
  wire net495;
  wire net496;
  wire net497;
  wire net498;
  wire net499;
  wire net500;
  wire net501;
  wire net502;
  wire net503;
  wire net504;
  wire net505;
  wire net506;
  wire net507;
  wire net508;
  wire net509;
  wire net510;
  wire net511;
  wire net512;
  wire net513;
  wire net514;
  wire net515;
  wire net516;
  wire net517;
  wire net518;
  wire net519;
  wire net520;
  wire net521;
  wire net522;
  wire net523;
  wire net524;
  wire net525;
  wire net526;
  wire net527;
  wire net528;
  wire net529;
  wire net530;
  wire net531;
  wire net532;
  wire net533;
  wire net534;
  wire net535;
  wire net536;
  wire net537;
  wire net538;
  wire net539;
  wire net540;
  wire net541;
  wire net542;
  wire net543;
  wire net544;
  wire net545;
  wire net546;
  wire net547;
  wire net548;
  wire net549;
  wire net550;

  assign uo_out[0] = net4;
  assign uo_out[1] = net5;
  assign uo_out[2] = net6;
  assign uo_out[3] = net7;
  assign uo_out[4] = net8;
  assign uo_out[5] = net9;
  assign uo_out[6] = net10;
  assign uo_out[7] = net11;
  assign uio_out[0] = 0;
  assign uio_oe[0] = 0;
  assign uio_out[1] = 0;
  assign uio_oe[1] = 0;
  assign uio_out[2] = 0;
  assign uio_oe[2] = 0;
  assign uio_out[3] = 0;
  assign uio_oe[3] = 0;
  assign uio_out[4] = 0;
  assign uio_oe[4] = 0;
  assign uio_out[5] = 0;
  assign uio_oe[5] = 0;
  assign uio_out[6] = 0;
  assign uio_oe[6] = 0;
  assign uio_out[7] = 0;
  assign uio_oe[7] = 0;

  mux_cell mux1 (
    .a (net17),
    .b (net2),
    .sel (net3),
    .out (net18)
  );
  dff_cell flipflop2 (
    .d (net19),
    .clk (net1),
    .q (net20),
    .notq (net21)
  );
  dff_cell flipflop3 (
    .d (net20),
    .clk (net1),
    .q (net22),
    .notq (net23)
  );
  dff_cell flipflop4 (
    .d (net22),
    .clk (net1),
    .q (net24),
    .notq (net25)
  );
  dff_cell flipflop5 (
    .d (net24),
    .clk (net1),
    .q (net26),
    .notq (net27)
  );
  dff_cell flipflop6 (
    .d (net26),
    .clk (net1),
    .q (net28),
    .notq (net29)
  );
  dff_cell flipflop7 (
    .d (net28),
    .clk (net1),
    .q (net30),
    .notq (net31)
  );
  dff_cell flipflop8 (
    .d (net30),
    .clk (net1),
    .q (net32),
    .notq (net33)
  );
  dff_cell flipflop9 (
    .d (net32),
    .clk (net1),
    .q (net34),
    .notq (net35)
  );
  dff_cell flipflop10 (
    .d (net34),
    .clk (net1),
    .q (net36),
    .notq (net37)
  );
  dff_cell flipflop11 (
    .d (net36),
    .clk (net1),
    .q (net38),
    .notq (net39)
  );
  dff_cell flipflop12 (
    .d (net38),
    .clk (net1),
    .q (net40),
    .notq (net41)
  );
  dff_cell flipflop13 (
    .d (net40),
    .clk (net1),
    .q (net42),
    .notq (net43)
  );
  dff_cell flipflop14 (
    .d (net42),
    .clk (net1),
    .q (net44),
    .notq (net45)
  );
  dff_cell flipflop15 (
    .d (net44),
    .clk (net1),
    .q (net46),
    .notq (net47)
  );
  dff_cell flipflop16 (
    .d (net46),
    .clk (net1),
    .q (net48),
    .notq (net49)
  );
  dff_cell flipflop1 (
    .d (net4),
    .clk (net1),
    .q (net19),
    .notq (net50)
  );
  or_cell gate1 (
    .a (net51),
    .b (net52),
    .out (net17)
  );
  and_cell gate2 (
    .a (net53),
    .b (net54),
    .out (net55)
  );
  and_cell gate4 (
    .a (net21),
    .b (net50),
    .out (net54)
  );
  and_cell gate5 (
    .a (net25),
    .b (net23),
    .out (net53)
  );
  and_cell gate6 (
    .a (net29),
    .b (net27),
    .out (net56)
  );
  and_cell gate9 (
    .a (net33),
    .b (net31),
    .out (net57)
  );
  and_cell gate10 (
    .a (net37),
    .b (net35),
    .out (net58)
  );
  and_cell gate11 (
    .a (net41),
    .b (net39),
    .out (net59)
  );
  and_cell gate12 (
    .a (net45),
    .b (net43),
    .out (net60)
  );
  and_cell gate13 (
    .a (net49),
    .b (net47),
    .out (net61)
  );
  and_cell gate14 (
    .a (net57),
    .b (net56),
    .out (net62)
  );
  and_cell gate15 (
    .a (net59),
    .b (net58),
    .out (net63)
  );
  and_cell gate16 (
    .a (net61),
    .b (net60),
    .out (net64)
  );
  and_cell gate17 (
    .a (net62),
    .b (net55),
    .out (net65)
  );
  and_cell gate19 (
    .a (net64),
    .b (net63),
    .out (net66)
  );
  and_cell gate20 (
    .a (net66),
    .b (net65),
    .out (net67)
  );
  dff_cell flipflop17 (
    .d (net48),
    .clk (net1),
    .q (net68),
    .notq (net69)
  );
  dff_cell flipflop18 (
    .d (net68),
    .clk (net1),
    .q (net70),
    .notq (net71)
  );
  dff_cell flipflop19 (
    .d (net70),
    .clk (net1),
    .q (net72),
    .notq (net73)
  );
  dff_cell flipflop20 (
    .d (net72),
    .clk (net1),
    .q (net74),
    .notq (net75)
  );
  dff_cell flipflop21 (
    .d (net74),
    .clk (net1),
    .q (net76),
    .notq (net77)
  );
  dff_cell flipflop22 (
    .d (net76),
    .clk (net1),
    .q (net78),
    .notq (net79)
  );
  dff_cell flipflop23 (
    .d (net78),
    .clk (net1),
    .q (net80),
    .notq (net81)
  );
  dff_cell flipflop24 (
    .d (net80),
    .clk (net1),
    .q (net82),
    .notq (net83)
  );
  dff_cell flipflop25 (
    .d (net82),
    .clk (net1),
    .q (net84),
    .notq (net85)
  );
  dff_cell flipflop26 (
    .d (net84),
    .clk (net1),
    .q (net86),
    .notq (net87)
  );
  dff_cell flipflop27 (
    .d (net86),
    .clk (net1),
    .q (net88),
    .notq (net89)
  );
  dff_cell flipflop28 (
    .d (net88),
    .clk (net1),
    .q (net90),
    .notq (net91)
  );
  dff_cell flipflop29 (
    .d (net90),
    .clk (net1),
    .q (net92),
    .notq (net93)
  );
  dff_cell flipflop30 (
    .d (net92),
    .clk (net1),
    .q (net94),
    .notq (net95)
  );
  dff_cell flipflop31 (
    .d (net94),
    .clk (net1),
    .q (net96),
    .notq (net97)
  );
  dff_cell flipflop32 (
    .d (net96),
    .clk (net1),
    .q (net98),
    .notq (net99)
  );
  and_cell gate23 (
    .a (net100),
    .b (net101),
    .out (net102)
  );
  and_cell gate24 (
    .a (net71),
    .b (net69),
    .out (net101)
  );
  and_cell gate25 (
    .a (net75),
    .b (net73),
    .out (net100)
  );
  and_cell gate26 (
    .a (net79),
    .b (net77),
    .out (net103)
  );
  and_cell gate32 (
    .a (net81),
    .b (net103),
    .out (net104)
  );
  and_cell gate35 (
    .a (net104),
    .b (net102),
    .out (net105)
  );
  and_cell gate37 (
    .a (net106),
    .b (net105),
    .out (net107)
  );
  and_cell and1 (
    .a (net107),
    .b (net67),
    .out (net108)
  );
  dff_cell flipflop33 (
    .d (net98),
    .clk (net1),
    .q (net109),
    .notq (net110)
  );
  dff_cell flipflop34 (
    .d (net109),
    .clk (net1),
    .q (net111),
    .notq (net112)
  );
  dff_cell flipflop35 (
    .d (net111),
    .clk (net1),
    .q (net113),
    .notq (net114)
  );
  dff_cell flipflop36 (
    .d (net113),
    .clk (net1),
    .q (net115),
    .notq (net116)
  );
  dff_cell flipflop37 (
    .d (net115),
    .clk (net1),
    .q (net117),
    .notq (net118)
  );
  dff_cell flipflop38 (
    .d (net117),
    .clk (net1),
    .q (net119),
    .notq (net120)
  );
  dff_cell flipflop39 (
    .d (net119),
    .clk (net1),
    .q (net121),
    .notq (net122)
  );
  dff_cell flipflop40 (
    .d (net121),
    .clk (net1),
    .q (net123),
    .notq (net124)
  );
  dff_cell flipflop41 (
    .d (net123),
    .clk (net1),
    .q (net125),
    .notq (net126)
  );
  dff_cell flipflop42 (
    .d (net125),
    .clk (net1),
    .q (net127),
    .notq (net128)
  );
  dff_cell flipflop43 (
    .d (net127),
    .clk (net1),
    .q (net129),
    .notq (net130)
  );
  dff_cell flipflop44 (
    .d (net129),
    .clk (net1),
    .q (net131),
    .notq (net132)
  );
  dff_cell flipflop45 (
    .d (net131),
    .clk (net1),
    .q (net133),
    .notq (net134)
  );
  dff_cell flipflop46 (
    .d (net133),
    .clk (net1),
    .q (net135),
    .notq (net136)
  );
  and_cell gate3 (
    .a (net137),
    .b (net138),
    .out (net139)
  );
  and_cell gate7 (
    .a (net85),
    .b (net83),
    .out (net138)
  );
  and_cell gate8 (
    .a (net89),
    .b (net87),
    .out (net137)
  );
  and_cell gate18 (
    .a (net93),
    .b (net91),
    .out (net140)
  );
  and_cell gate21 (
    .a (net97),
    .b (net95),
    .out (net141)
  );
  and_cell gate22 (
    .a (net110),
    .b (net99),
    .out (net142)
  );
  and_cell gate27 (
    .a (net114),
    .b (net112),
    .out (net143)
  );
  and_cell gate28 (
    .a (net118),
    .b (net116),
    .out (net144)
  );
  and_cell gate29 (
    .a (net122),
    .b (net120),
    .out (net145)
  );
  and_cell gate30 (
    .a (net141),
    .b (net140),
    .out (net146)
  );
  and_cell gate31 (
    .a (net143),
    .b (net142),
    .out (net147)
  );
  and_cell gate33 (
    .a (net145),
    .b (net144),
    .out (net148)
  );
  and_cell gate34 (
    .a (net146),
    .b (net139),
    .out (net149)
  );
  and_cell gate36 (
    .a (net148),
    .b (net147),
    .out (net150)
  );
  and_cell gate38 (
    .a (net150),
    .b (net149),
    .out (net151)
  );
  and_cell gate39 (
    .a (net152),
    .b (net153),
    .out (net154)
  );
  and_cell gate40 (
    .a (net126),
    .b (net124),
    .out (net153)
  );
  and_cell gate41 (
    .a (net130),
    .b (net128),
    .out (net152)
  );
  and_cell gate42 (
    .a (net134),
    .b (net132),
    .out (net155)
  );
  and_cell gate43 (
    .a (net136),
    .b (net155),
    .out (net156)
  );
  and_cell gate44 (
    .a (net156),
    .b (net154),
    .out (net106)
  );
  and_cell gate45 (
    .a (net157),
    .b (net151),
    .out (net158)
  );
  dff_cell flipflop47 (
    .d (net135),
    .clk (net1),
    .q (net159),
    .notq (net160)
  );
  dff_cell flipflop48 (
    .d (net159),
    .clk (net1),
    .q (net161),
    .notq (net162)
  );
  dff_cell flipflop49 (
    .d (net161),
    .clk (net1),
    .q (net163),
    .notq (net164)
  );
  dff_cell flipflop50 (
    .d (net163),
    .clk (net1),
    .q (net165),
    .notq (net166)
  );
  dff_cell flipflop51 (
    .d (net165),
    .clk (net1),
    .q (net167),
    .notq (net168)
  );
  dff_cell flipflop52 (
    .d (net167),
    .clk (net1),
    .q (net169),
    .notq (net170)
  );
  dff_cell flipflop53 (
    .d (net169),
    .clk (net1),
    .q (net171),
    .notq (net172)
  );
  dff_cell flipflop54 (
    .d (net171),
    .clk (net1),
    .q (net173),
    .notq (net174)
  );
  dff_cell flipflop55 (
    .d (net173),
    .clk (net1),
    .q (net175),
    .notq (net176)
  );
  dff_cell flipflop56 (
    .d (net175),
    .clk (net1),
    .q (net177),
    .notq (net178)
  );
  dff_cell flipflop57 (
    .d (net177),
    .clk (net1),
    .q (net179),
    .notq (net180)
  );
  dff_cell flipflop58 (
    .d (net179),
    .clk (net1),
    .q (net181),
    .notq (net182)
  );
  dff_cell flipflop59 (
    .d (net181),
    .clk (net1),
    .q (net183),
    .notq (net184)
  );
  dff_cell flipflop60 (
    .d (net183),
    .clk (net1),
    .q (net185),
    .notq (net186)
  );
  dff_cell flipflop61 (
    .d (net185),
    .clk (net1),
    .q (net187),
    .notq (net188)
  );
  dff_cell flipflop62 (
    .d (net187),
    .clk (net1),
    .q (net189),
    .notq (net190)
  );
  and_cell gate46 (
    .a (net191),
    .b (net192),
    .out (net193)
  );
  and_cell gate47 (
    .a (net162),
    .b (net160),
    .out (net192)
  );
  and_cell gate48 (
    .a (net166),
    .b (net164),
    .out (net191)
  );
  and_cell gate49 (
    .a (net170),
    .b (net168),
    .out (net194)
  );
  and_cell gate50 (
    .a (net174),
    .b (net172),
    .out (net195)
  );
  and_cell gate51 (
    .a (net178),
    .b (net176),
    .out (net196)
  );
  and_cell gate52 (
    .a (net182),
    .b (net180),
    .out (net197)
  );
  and_cell gate53 (
    .a (net186),
    .b (net184),
    .out (net198)
  );
  and_cell gate54 (
    .a (net190),
    .b (net188),
    .out (net199)
  );
  and_cell gate55 (
    .a (net195),
    .b (net194),
    .out (net200)
  );
  and_cell gate56 (
    .a (net197),
    .b (net196),
    .out (net201)
  );
  and_cell gate57 (
    .a (net199),
    .b (net198),
    .out (net202)
  );
  and_cell gate58 (
    .a (net200),
    .b (net193),
    .out (net203)
  );
  and_cell gate59 (
    .a (net202),
    .b (net201),
    .out (net204)
  );
  and_cell gate60 (
    .a (net204),
    .b (net203),
    .out (net157)
  );
  dff_cell flipflop63 (
    .d (net189),
    .clk (net1),
    .q (net205),
    .notq (net206)
  );
  dff_cell flipflop64 (
    .d (net205),
    .clk (net1),
    .q (net207),
    .notq (net208)
  );
  dff_cell flipflop65 (
    .d (net207),
    .clk (net1),
    .q (net7),
    .notq (net209)
  );
  dff_cell flipflop66 (
    .d (net7),
    .clk (net1),
    .q (net210),
    .notq (net211)
  );
  dff_cell flipflop67 (
    .d (net210),
    .clk (net1),
    .q (net212),
    .notq (net213)
  );
  dff_cell flipflop68 (
    .d (net212),
    .clk (net1),
    .q (net5),
    .notq (net214)
  );
  dff_cell flipflop69 (
    .d (net5),
    .clk (net1),
    .q (net215),
    .notq (net216)
  );
  dff_cell flipflop70 (
    .d (net215),
    .clk (net1),
    .q (net217),
    .notq (net218)
  );
  dff_cell flipflop71 (
    .d (net217),
    .clk (net1),
    .q (net219),
    .notq (net220)
  );
  dff_cell flipflop72 (
    .d (net219),
    .clk (net1),
    .q (net221),
    .notq (net222)
  );
  dff_cell flipflop73 (
    .d (net221),
    .clk (net1),
    .q (net223),
    .notq (net224)
  );
  dff_cell flipflop74 (
    .d (net223),
    .clk (net1),
    .q (net225),
    .notq (net226)
  );
  dff_cell flipflop75 (
    .d (net225),
    .clk (net1),
    .q (net227),
    .notq (net228)
  );
  dff_cell flipflop76 (
    .d (net227),
    .clk (net1),
    .q (net229),
    .notq (net230)
  );
  dff_cell flipflop77 (
    .d (net229),
    .clk (net1),
    .q (net231),
    .notq (net232)
  );
  dff_cell flipflop78 (
    .d (net231),
    .clk (net1),
    .q (net233),
    .notq (net234)
  );
  and_cell gate61 (
    .a (net235),
    .b (net236),
    .out (net237)
  );
  and_cell gate62 (
    .a (net208),
    .b (net206),
    .out (net236)
  );
  and_cell gate63 (
    .a (net211),
    .b (net209),
    .out (net235)
  );
  and_cell gate64 (
    .a (net214),
    .b (net213),
    .out (net238)
  );
  and_cell gate65 (
    .a (net216),
    .b (net238),
    .out (net239)
  );
  and_cell gate66 (
    .a (net239),
    .b (net237),
    .out (net240)
  );
  and_cell gate67 (
    .a (net241),
    .b (net240),
    .out (net242)
  );
  and_cell and2 (
    .a (net243),
    .b (net242),
    .out (net244)
  );
  dff_cell flipflop79 (
    .d (net233),
    .clk (net1),
    .q (net245),
    .notq (net246)
  );
  dff_cell flipflop80 (
    .d (net245),
    .clk (net1),
    .q (net247),
    .notq (net248)
  );
  dff_cell flipflop81 (
    .d (net247),
    .clk (net1),
    .q (net249),
    .notq (net250)
  );
  dff_cell flipflop82 (
    .d (net249),
    .clk (net1),
    .q (net251),
    .notq (net252)
  );
  dff_cell flipflop83 (
    .d (net251),
    .clk (net1),
    .q (net253),
    .notq (net254)
  );
  dff_cell flipflop84 (
    .d (net253),
    .clk (net1),
    .q (net255),
    .notq (net256)
  );
  dff_cell flipflop85 (
    .d (net255),
    .clk (net1),
    .q (net257),
    .notq (net258)
  );
  dff_cell flipflop86 (
    .d (net257),
    .clk (net1),
    .q (net259),
    .notq (net260)
  );
  dff_cell flipflop87 (
    .d (net259),
    .clk (net1),
    .q (net261),
    .notq (net262)
  );
  dff_cell flipflop88 (
    .d (net261),
    .clk (net1),
    .q (net263),
    .notq (net264)
  );
  dff_cell flipflop89 (
    .d (net263),
    .clk (net1),
    .q (net265),
    .notq (net266)
  );
  dff_cell flipflop90 (
    .d (net265),
    .clk (net1),
    .q (net267),
    .notq (net268)
  );
  dff_cell flipflop91 (
    .d (net267),
    .clk (net1),
    .q (net269),
    .notq (net270)
  );
  dff_cell flipflop92 (
    .d (net269),
    .clk (net1),
    .q (net8),
    .notq (net271)
  );
  and_cell gate68 (
    .a (net272),
    .b (net273),
    .out (net274)
  );
  and_cell gate69 (
    .a (net220),
    .b (net218),
    .out (net273)
  );
  and_cell gate70 (
    .a (net224),
    .b (net222),
    .out (net272)
  );
  and_cell gate71 (
    .a (net228),
    .b (net226),
    .out (net275)
  );
  and_cell gate72 (
    .a (net232),
    .b (net230),
    .out (net276)
  );
  and_cell gate73 (
    .a (net246),
    .b (net234),
    .out (net277)
  );
  and_cell gate74 (
    .a (net250),
    .b (net248),
    .out (net278)
  );
  and_cell gate75 (
    .a (net254),
    .b (net252),
    .out (net279)
  );
  and_cell gate76 (
    .a (net258),
    .b (net256),
    .out (net280)
  );
  and_cell gate77 (
    .a (net276),
    .b (net275),
    .out (net281)
  );
  and_cell gate78 (
    .a (net278),
    .b (net277),
    .out (net282)
  );
  and_cell gate79 (
    .a (net280),
    .b (net279),
    .out (net283)
  );
  and_cell gate80 (
    .a (net281),
    .b (net274),
    .out (net284)
  );
  and_cell gate81 (
    .a (net283),
    .b (net282),
    .out (net285)
  );
  and_cell gate82 (
    .a (net285),
    .b (net284),
    .out (net243)
  );
  and_cell gate83 (
    .a (net286),
    .b (net287),
    .out (net288)
  );
  and_cell gate84 (
    .a (net262),
    .b (net260),
    .out (net287)
  );
  and_cell gate85 (
    .a (net266),
    .b (net264),
    .out (net286)
  );
  and_cell gate86 (
    .a (net270),
    .b (net268),
    .out (net289)
  );
  and_cell gate87 (
    .a (net271),
    .b (net289),
    .out (net290)
  );
  and_cell gate88 (
    .a (net290),
    .b (net288),
    .out (net241)
  );
  and_cell and3 (
    .a (net244),
    .b (net158),
    .out (net291)
  );
  and_cell and4 (
    .a (net291),
    .b (net108),
    .out (net292)
  );
  dff_cell flipflop93 (
    .d (net293),
    .clk (net1),
    .q (net294),
    .notq (net295)
  );
  dff_cell flipflop94 (
    .d (net294),
    .clk (net1),
    .q (net296),
    .notq (net297)
  );
  dff_cell flipflop95 (
    .d (net296),
    .clk (net1),
    .q (net298),
    .notq (net299)
  );
  dff_cell flipflop96 (
    .d (net298),
    .clk (net1),
    .q (net300),
    .notq (net301)
  );
  dff_cell flipflop97 (
    .d (net300),
    .clk (net1),
    .q (net302),
    .notq (net303)
  );
  dff_cell flipflop98 (
    .d (net302),
    .clk (net1),
    .q (net304),
    .notq (net305)
  );
  dff_cell flipflop99 (
    .d (net304),
    .clk (net1),
    .q (net306),
    .notq (net307)
  );
  dff_cell flipflop100 (
    .d (net306),
    .clk (net1),
    .q (net308),
    .notq (net309)
  );
  dff_cell flipflop101 (
    .d (net308),
    .clk (net1),
    .q (net310),
    .notq (net311)
  );
  and_cell gate89 (
    .a (net312),
    .b (net313),
    .out (net314)
  );
  dff_cell flipflop102 (
    .d (net310),
    .clk (net1),
    .q (net315),
    .notq (net316)
  );
  dff_cell flipflop103 (
    .d (net315),
    .clk (net1),
    .q (net317),
    .notq (net318)
  );
  dff_cell flipflop104 (
    .d (net317),
    .clk (net1),
    .q (net319),
    .notq (net320)
  );
  dff_cell flipflop105 (
    .d (net319),
    .clk (net1),
    .q (net321),
    .notq (net322)
  );
  dff_cell flipflop106 (
    .d (net321),
    .clk (net1),
    .q (net323),
    .notq (net324)
  );
  dff_cell flipflop107 (
    .d (net323),
    .clk (net1),
    .q (net325),
    .notq (net326)
  );
  dff_cell flipflop108 (
    .d (net325),
    .clk (net1),
    .q (net327),
    .notq (net328)
  );
  dff_cell flipflop109 (
    .d (net327),
    .clk (net1),
    .q (net329),
    .notq (net330)
  );
  dff_cell flipflop110 (
    .d (net329),
    .clk (net1),
    .q (net331),
    .notq (net332)
  );
  dff_cell flipflop111 (
    .d (net331),
    .clk (net1),
    .q (net333),
    .notq (net334)
  );
  dff_cell flipflop112 (
    .d (net333),
    .clk (net1),
    .q (net335),
    .notq (net336)
  );
  dff_cell flipflop113 (
    .d (net335),
    .clk (net1),
    .q (net337),
    .notq (net338)
  );
  and_cell gate90 (
    .a (net339),
    .b (net340),
    .out (net341)
  );
  and_cell gate91 (
    .a (net297),
    .b (net295),
    .out (net340)
  );
  and_cell gate92 (
    .a (net301),
    .b (net299),
    .out (net339)
  );
  and_cell gate93 (
    .a (net305),
    .b (net303),
    .out (net342)
  );
  and_cell gate94 (
    .a (net309),
    .b (net307),
    .out (net343)
  );
  and_cell gate95 (
    .a (net316),
    .b (net311),
    .out (net344)
  );
  and_cell gate96 (
    .a (net320),
    .b (net318),
    .out (net345)
  );
  and_cell gate97 (
    .a (net324),
    .b (net322),
    .out (net346)
  );
  and_cell gate98 (
    .a (net328),
    .b (net326),
    .out (net347)
  );
  and_cell gate99 (
    .a (net343),
    .b (net342),
    .out (net348)
  );
  and_cell gate100 (
    .a (net345),
    .b (net344),
    .out (net349)
  );
  and_cell gate101 (
    .a (net347),
    .b (net346),
    .out (net350)
  );
  and_cell gate102 (
    .a (net348),
    .b (net341),
    .out (net351)
  );
  and_cell gate103 (
    .a (net350),
    .b (net349),
    .out (net352)
  );
  and_cell gate104 (
    .a (net352),
    .b (net351),
    .out (net353)
  );
  and_cell gate105 (
    .a (net354),
    .b (net355),
    .out (net356)
  );
  and_cell gate106 (
    .a (net332),
    .b (net330),
    .out (net355)
  );
  and_cell gate107 (
    .a (net336),
    .b (net334),
    .out (net354)
  );
  and_cell gate110 (
    .a (net338),
    .b (net356),
    .out (net313)
  );
  dff_cell flipflop114 (
    .d (net337),
    .clk (net1),
    .q (net357),
    .notq (net358)
  );
  dff_cell flipflop115 (
    .d (net357),
    .clk (net1),
    .q (net359),
    .notq (net360)
  );
  dff_cell flipflop116 (
    .d (net359),
    .clk (net1),
    .q (net361),
    .notq (net362)
  );
  dff_cell flipflop117 (
    .d (net361),
    .clk (net1),
    .q (net363),
    .notq (net364)
  );
  dff_cell flipflop118 (
    .d (net363),
    .clk (net1),
    .q (net365),
    .notq (net366)
  );
  dff_cell flipflop119 (
    .d (net365),
    .clk (net1),
    .q (net367),
    .notq (net368)
  );
  dff_cell flipflop120 (
    .d (net367),
    .clk (net1),
    .q (net369),
    .notq (net370)
  );
  dff_cell flipflop121 (
    .d (net369),
    .clk (net1),
    .q (net371),
    .notq (net372)
  );
  dff_cell flipflop122 (
    .d (net371),
    .clk (net1),
    .q (net373),
    .notq (net374)
  );
  dff_cell flipflop123 (
    .d (net373),
    .clk (net1),
    .q (net375),
    .notq (net376)
  );
  dff_cell flipflop124 (
    .d (net375),
    .clk (net1),
    .q (net377),
    .notq (net378)
  );
  dff_cell flipflop125 (
    .d (net377),
    .clk (net1),
    .q (net379),
    .notq (net380)
  );
  dff_cell flipflop126 (
    .d (net379),
    .clk (net1),
    .q (net381),
    .notq (net382)
  );
  dff_cell flipflop127 (
    .d (net381),
    .clk (net1),
    .q (net383),
    .notq (net384)
  );
  dff_cell flipflop128 (
    .d (net383),
    .clk (net1),
    .q (net385),
    .notq (net386)
  );
  dff_cell flipflop129 (
    .d (net385),
    .clk (net1),
    .q (net387),
    .notq (net388)
  );
  dff_cell flipflop130 (
    .d (net387),
    .clk (net1),
    .q (net389),
    .notq (net390)
  );
  dff_cell flipflop131 (
    .d (net389),
    .clk (net1),
    .q (net391),
    .notq (net392)
  );
  dff_cell flipflop132 (
    .d (net391),
    .clk (net1),
    .q (net393),
    .notq (net394)
  );
  dff_cell flipflop133 (
    .d (net393),
    .clk (net1),
    .q (net395),
    .notq (net396)
  );
  dff_cell flipflop134 (
    .d (net395),
    .clk (net1),
    .q (net397),
    .notq (net398)
  );
  and_cell gate109 (
    .a (net399),
    .b (net400),
    .out (net401)
  );
  and_cell gate111 (
    .a (net360),
    .b (net358),
    .out (net400)
  );
  and_cell gate112 (
    .a (net364),
    .b (net362),
    .out (net399)
  );
  and_cell gate113 (
    .a (net368),
    .b (net366),
    .out (net402)
  );
  and_cell gate114 (
    .a (net372),
    .b (net370),
    .out (net403)
  );
  and_cell gate115 (
    .a (net376),
    .b (net374),
    .out (net404)
  );
  and_cell gate116 (
    .a (net380),
    .b (net378),
    .out (net405)
  );
  and_cell gate117 (
    .a (net384),
    .b (net382),
    .out (net406)
  );
  and_cell gate118 (
    .a (net388),
    .b (net386),
    .out (net407)
  );
  and_cell gate119 (
    .a (net403),
    .b (net402),
    .out (net408)
  );
  and_cell gate120 (
    .a (net405),
    .b (net404),
    .out (net409)
  );
  and_cell gate121 (
    .a (net407),
    .b (net406),
    .out (net410)
  );
  and_cell gate122 (
    .a (net408),
    .b (net401),
    .out (net411)
  );
  and_cell gate123 (
    .a (net410),
    .b (net409),
    .out (net412)
  );
  and_cell gate124 (
    .a (net412),
    .b (net411),
    .out (net413)
  );
  and_cell gate125 (
    .a (net414),
    .b (net415),
    .out (net416)
  );
  and_cell gate126 (
    .a (net392),
    .b (net390),
    .out (net415)
  );
  and_cell gate127 (
    .a (net396),
    .b (net394),
    .out (net414)
  );
  and_cell gate128 (
    .a (net398),
    .b (net416),
    .out (net312)
  );
  dff_cell flipflop135 (
    .d (net397),
    .clk (net1),
    .q (net417),
    .notq (net418)
  );
  dff_cell flipflop136 (
    .d (net417),
    .clk (net1),
    .q (net419),
    .notq (net420)
  );
  dff_cell flipflop137 (
    .d (net419),
    .clk (net1),
    .q (net421),
    .notq (net422)
  );
  dff_cell flipflop138 (
    .d (net421),
    .clk (net1),
    .q (net423),
    .notq (net424)
  );
  dff_cell flipflop139 (
    .d (net423),
    .clk (net1),
    .q (net425),
    .notq (net426)
  );
  dff_cell flipflop140 (
    .d (net425),
    .clk (net1),
    .q (net427),
    .notq (net428)
  );
  dff_cell flipflop141 (
    .d (net427),
    .clk (net1),
    .q (net429),
    .notq (net430)
  );
  dff_cell flipflop142 (
    .d (net429),
    .clk (net1),
    .q (net431),
    .notq (net432)
  );
  dff_cell flipflop143 (
    .d (net431),
    .clk (net1),
    .q (net433),
    .notq (net434)
  );
  and_cell gate108 (
    .a (net435),
    .b (net436),
    .out (net437)
  );
  dff_cell flipflop144 (
    .d (net433),
    .clk (net1),
    .q (net438),
    .notq (net439)
  );
  dff_cell flipflop145 (
    .d (net438),
    .clk (net1),
    .q (net440),
    .notq (net441)
  );
  dff_cell flipflop146 (
    .d (net440),
    .clk (net1),
    .q (net442),
    .notq (net443)
  );
  dff_cell flipflop147 (
    .d (net442),
    .clk (net1),
    .q (net444),
    .notq (net445)
  );
  dff_cell flipflop148 (
    .d (net444),
    .clk (net1),
    .q (net446),
    .notq (net447)
  );
  dff_cell flipflop149 (
    .d (net446),
    .clk (net1),
    .q (net448),
    .notq (net449)
  );
  dff_cell flipflop150 (
    .d (net448),
    .clk (net1),
    .q (net450),
    .notq (net451)
  );
  dff_cell flipflop151 (
    .d (net450),
    .clk (net1),
    .q (net452),
    .notq (net453)
  );
  dff_cell flipflop152 (
    .d (net452),
    .clk (net1),
    .q (net454),
    .notq (net455)
  );
  dff_cell flipflop153 (
    .d (net454),
    .clk (net1),
    .q (net456),
    .notq (net457)
  );
  dff_cell flipflop154 (
    .d (net456),
    .clk (net1),
    .q (net458),
    .notq (net459)
  );
  dff_cell flipflop155 (
    .d (net458),
    .clk (net1),
    .q (net460),
    .notq (net461)
  );
  and_cell gate129 (
    .a (net462),
    .b (net463),
    .out (net464)
  );
  and_cell gate130 (
    .a (net420),
    .b (net418),
    .out (net463)
  );
  and_cell gate131 (
    .a (net424),
    .b (net422),
    .out (net462)
  );
  and_cell gate132 (
    .a (net428),
    .b (net426),
    .out (net465)
  );
  and_cell gate133 (
    .a (net432),
    .b (net430),
    .out (net466)
  );
  and_cell gate134 (
    .a (net439),
    .b (net434),
    .out (net467)
  );
  and_cell gate135 (
    .a (net443),
    .b (net441),
    .out (net468)
  );
  and_cell gate136 (
    .a (net447),
    .b (net445),
    .out (net469)
  );
  and_cell gate137 (
    .a (net451),
    .b (net449),
    .out (net470)
  );
  and_cell gate138 (
    .a (net466),
    .b (net465),
    .out (net471)
  );
  and_cell gate139 (
    .a (net468),
    .b (net467),
    .out (net472)
  );
  and_cell gate140 (
    .a (net470),
    .b (net469),
    .out (net473)
  );
  and_cell gate141 (
    .a (net471),
    .b (net464),
    .out (net474)
  );
  and_cell gate142 (
    .a (net473),
    .b (net472),
    .out (net475)
  );
  and_cell gate143 (
    .a (net475),
    .b (net474),
    .out (net476)
  );
  and_cell gate144 (
    .a (net477),
    .b (net478),
    .out (net479)
  );
  and_cell gate145 (
    .a (net455),
    .b (net453),
    .out (net478)
  );
  and_cell gate146 (
    .a (net459),
    .b (net457),
    .out (net477)
  );
  and_cell gate147 (
    .a (net461),
    .b (net479),
    .out (net436)
  );
  dff_cell flipflop156 (
    .d (net460),
    .clk (net1),
    .q (net480),
    .notq (net481)
  );
  dff_cell flipflop157 (
    .d (net480),
    .clk (net1),
    .q (net482),
    .notq (net483)
  );
  dff_cell flipflop158 (
    .d (net482),
    .clk (net1),
    .q (net484),
    .notq (net485)
  );
  dff_cell flipflop159 (
    .d (net484),
    .clk (net1),
    .q (net486),
    .notq (net487)
  );
  dff_cell flipflop160 (
    .d (net486),
    .clk (net1),
    .q (net488),
    .notq (net489)
  );
  dff_cell flipflop161 (
    .d (net488),
    .clk (net1),
    .q (net9),
    .notq (net490)
  );
  dff_cell flipflop162 (
    .d (net9),
    .clk (net1),
    .q (net491),
    .notq (net492)
  );
  dff_cell flipflop163 (
    .d (net491),
    .clk (net1),
    .q (net493),
    .notq (net494)
  );
  dff_cell flipflop164 (
    .d (net493),
    .clk (net1),
    .q (net495),
    .notq (net496)
  );
  dff_cell flipflop165 (
    .d (net495),
    .clk (net1),
    .q (net497),
    .notq (net498)
  );
  dff_cell flipflop166 (
    .d (net497),
    .clk (net1),
    .q (net499),
    .notq (net500)
  );
  dff_cell flipflop167 (
    .d (net499),
    .clk (net1),
    .q (net501),
    .notq (net502)
  );
  dff_cell flipflop168 (
    .d (net501),
    .clk (net1),
    .q (net503),
    .notq (net504)
  );
  dff_cell flipflop169 (
    .d (net503),
    .clk (net1),
    .q (net505),
    .notq (net506)
  );
  dff_cell flipflop170 (
    .d (net505),
    .clk (net1),
    .q (net507),
    .notq (net508)
  );
  dff_cell flipflop171 (
    .d (net507),
    .clk (net1),
    .q (net509),
    .notq (net510)
  );
  dff_cell flipflop172 (
    .d (net509),
    .clk (net1),
    .q (net511),
    .notq (net512)
  );
  dff_cell flipflop173 (
    .d (net511),
    .clk (net1),
    .q (net513),
    .notq (net514)
  );
  dff_cell flipflop174 (
    .d (net513),
    .clk (net1),
    .q (net515),
    .notq (net516)
  );
  dff_cell flipflop175 (
    .d (net515),
    .clk (net1),
    .q (net517),
    .notq (net518)
  );
  dff_cell flipflop176 (
    .d (net517),
    .clk (net1),
    .q (net10),
    .notq (net519)
  );
  and_cell gate148 (
    .a (net520),
    .b (net521),
    .out (net522)
  );
  and_cell gate149 (
    .a (net483),
    .b (net481),
    .out (net521)
  );
  and_cell gate150 (
    .a (net487),
    .b (net485),
    .out (net520)
  );
  and_cell gate151 (
    .a (net490),
    .b (net489),
    .out (net523)
  );
  and_cell gate152 (
    .a (net494),
    .b (net492),
    .out (net524)
  );
  and_cell gate153 (
    .a (net498),
    .b (net496),
    .out (net525)
  );
  and_cell gate154 (
    .a (net502),
    .b (net500),
    .out (net526)
  );
  and_cell gate155 (
    .a (net506),
    .b (net504),
    .out (net527)
  );
  and_cell gate156 (
    .a (net510),
    .b (net508),
    .out (net528)
  );
  and_cell gate157 (
    .a (net524),
    .b (net523),
    .out (net529)
  );
  and_cell gate158 (
    .a (net526),
    .b (net525),
    .out (net530)
  );
  and_cell gate159 (
    .a (net528),
    .b (net527),
    .out (net531)
  );
  and_cell gate160 (
    .a (net529),
    .b (net522),
    .out (net532)
  );
  and_cell gate161 (
    .a (net531),
    .b (net530),
    .out (net533)
  );
  and_cell gate162 (
    .a (net533),
    .b (net532),
    .out (net534)
  );
  and_cell gate163 (
    .a (net535),
    .b (net536),
    .out (net537)
  );
  and_cell gate164 (
    .a (net514),
    .b (net512),
    .out (net536)
  );
  and_cell gate165 (
    .a (net518),
    .b (net516),
    .out (net535)
  );
  and_cell gate166 (
    .a (net519),
    .b (net537),
    .out (net435)
  );
  and_cell gate167 (
    .a (net314),
    .b (net353),
    .out (net538)
  );
  and_cell gate168 (
    .a (net413),
    .b (net538),
    .out (net539)
  );
  and_cell gate169 (
    .a (net437),
    .b (net476),
    .out (net540)
  );
  and_cell gate170 (
    .a (net534),
    .b (net540),
    .out (net541)
  );
  and_cell gate171 (
    .a (net541),
    .b (net539),
    .out (net542)
  );
  and_cell gate172 (
    .a (net542),
    .b (net292),
    .out (net543)
  );
  dff_cell flipflop0 (
    .d (net18),
    .clk (net1),
    .q (net4),
    .notq (net544)
  );
  and_cell gate173 (
    .a (net543),
    .b (net544),
    .out (net51)
  );
  and_cell and5 (
    .a (net267),
    .b (net269),
    .out (net545)
  );
  xor_cell xor1 (
    .a (net8),
    .b (net7),
    .out (net546)
  );
  xor_cell xor2 (
    .a (net546),
    .b (net545),
    .out (net547)
  );
  xor_cell xor3 (
    .a (net507),
    .b (net547),
    .out (net548)
  );
  mux_cell mux2 (
    .a (net548),
    .b (net8),
    .sel (net3),
    .out (net293)
  );
  and_cell and6 (
    .a (net515),
    .b (net517),
    .out (net549)
  );
  xor_cell xor4 (
    .a (net10),
    .b (net9),
    .out (net550)
  );
  xor_cell xor5 (
    .a (net550),
    .b (net549),
    .out (net6)
  );
  xor_cell xor6 (
    .a (net550),
    .b (net546),
    .out (net11)
  );
  xor_cell xor7 (
    .a (net6),
    .b (net5),
    .out (net52)
  );
endmodule
